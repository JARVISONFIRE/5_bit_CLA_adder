* SPICE3 file created from DFF.ext - technology: scmos

.option scale=90n

M1000 out a_131_26# vdd w_156_21# pfet w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1001 stage_2_out stage_1_out a_93_9# Gnd nfet w=4 l=2
+  ad=20p pd=18u as=12p ps=10u
M1002 a_131_9# stage_2_out gnd Gnd nfet w=4 l=2
+  ad=12p pd=10u as=20p ps=18u
M1003 out a_131_26# gnd Gnd nfet w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1004 a_50_26# D vdd w_37_20# pfet w=8 l=2
+  ad=24p pd=14u as=40p ps=26u
M1005 a_131_26# stage_2_out vdd w_118_20# pfet w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1006 a_93_9# clk gnd Gnd nfet w=4 l=2
+  ad=12p pd=10u as=20p ps=18u
M1007 stage_2_out clk vdd w_80_20# pfet w=8 l=2
+  ad=40p pd=26u as=40p ps=26u
M1008 stage_1_out D gnd Gnd nfet w=4 l=2
+  ad=20p pd=18u as=20p ps=18u
M1009 a_131_26# clk a_131_9# Gnd nfet w=4 l=2
+  ad=20p pd=18u as=12p ps=10u
M1010 stage_1_out clk a_50_26# w_37_20# pfet w=8 l=2
+  ad=40p pd=26u as=24p ps=14u
C0 gnd a_93_9# 0.07426f
C1 w_37_20# D 0.02417f
C2 clk a_131_26# 0.17427f
C3 D vdd 0.03468f
C4 out w_156_21# 0.00935f
C5 gnd a_131_9# 0.08252f
C6 w_37_20# clk 0.03952f
C7 clk vdd 0.18083f
C8 stage_1_out clk 0.10999f
C9 stage_2_out vdd 0.13531f
C10 stage_1_out stage_2_out 0.15132f
C11 gnd D 0.04309f
C12 a_131_26# vdd 0.12809f
C13 a_50_26# vdd 0.10605f
C14 gnd clk 0.05789f
C15 a_50_26# stage_1_out 0.08248f
C16 w_37_20# vdd 0.00842f
C17 w_37_20# stage_1_out 0.00794f
C18 w_80_20# clk 0.02124f
C19 stage_1_out vdd 0.02357f
C20 out a_131_26# 0.0591f
C21 gnd stage_2_out 0.09001f
C22 w_118_20# clk 0
C23 w_80_20# stage_2_out 0.01186f
C24 out vdd 0.12374f
C25 a_93_9# stage_2_out 0.04124f
C26 gnd a_131_26# 0.09794f
C27 w_118_20# stage_2_out 0.02507f
C28 w_156_21# clk 0
C29 stage_1_out gnd 0.32172f
C30 w_118_20# a_131_26# 0.01186f
C31 w_80_20# vdd 0.00839f
C32 D clk 0.02644f
C33 a_131_9# a_131_26# 0.04124f
C34 stage_1_out w_80_20# 0
C35 stage_1_out a_93_9# 0.00603f
C36 out gnd 0.0825f
C37 w_156_21# a_131_26# 0.02707f
C38 w_118_20# vdd 0.00841f
C39 w_156_21# vdd 0.03739f
C40 clk stage_2_out 0.03022f
C41 a_131_9# 0 0.0042f **FLOATING
C42 a_93_9# 0 0.00422f **FLOATING
C43 gnd 0 0.52109f **FLOATING
C44 out 0 0.07734f **FLOATING
C45 stage_1_out 0 0.66306f **FLOATING
C46 a_50_26# 0 0.00438f **FLOATING
C47 vdd 0 0.50064f **FLOATING
C48 a_131_26# 0 0.28752f **FLOATING
C49 stage_2_out 0 0.25774f **FLOATING
C50 clk 0 1.85008f **FLOATING
C51 D 0 0.14714f **FLOATING
C52 w_156_21# 0 0.57753f **FLOATING
C53 w_118_20# 0 0.48211f **FLOATING
C54 w_80_20# 0 0.48211f **FLOATING
C55 w_37_20# 0 0.64282f **FLOATING
