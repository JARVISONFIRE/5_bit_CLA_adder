* =========================================================
* CPL XOR + DOMINO CLA - 180nm - Comparison Testbench
* Save as: CPL_XOR_domino_comparison.cir
* =========================================================
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.09u
.param WN = {4*LAMBDA}
.param WP = {8*LAMBDA}
.global gnd

* --- Supplies & Stimuli (same as CMOS file) ---
Vdd vdd 0 'SUPPLY'
Va2 a2 0 PULSE(0 'SUPPLY' 25n 100p 100p 10n 20n)
Vb2 b2 0 PULSE(0 'SUPPLY' 35n 100p 100p 20n 40n)
Va1 a1 0 PULSE(0 'SUPPLY' 25n 100p 100p 5n 10n)
Vb1 b1 0 PULSE(0 'SUPPLY' 30n 100p 100p 10n 20n)
Va0 a0 0 PULSE(0 'SUPPLY' 25n 100p 100p 2.5n 5n)
Vb0 b0 0 PULSE(0 'SUPPLY' 27.5n 100p 100p 5n 10n)
Vcin c0 0 PULSE(0 'SUPPLY' 55n 100p 100p 10n 20n)
Vclk clk 0 PULSE(0 'SUPPLY' 0 100p 100p 10n 20n)

* --- Basic CMOS inverter (buffers) ---
.subckt CMOS_INV A Y vdd gnd
Mpi Y A vdd vdd CMOSP W={WP} L={2*LAMBDA}
Mni Y A gnd gnd CMOSN W={WN} L={2*LAMBDA}
.ends

* --- CPL XOR (pass-transistor style) with level-restoring buffer
* Note: We generate complements via inverters locally for robustness
.subckt CPL_XOR2 A B Y vdd gnd
* generate complements
Xainv A A_n vdd gnd CMOS_INV
Xbinv B B_n vdd gnd CMOS_INV

* pass-transistor tree (simple 4T-ish implementation) producing xint
Mpx1 xint B A_n 0 0 CMOSN W={WN} L={2*LAMBDA}
Mpx2 xint B_n A 0 0 CMOSN W={WN} L={2*LAMBDA}
* level-restoring buffer to full swing
Xbuf_x xint Y vdd gnd CMOS_INV
.ends

* --- CPL AND (pass-transistor + buffer) producing G
.subckt CPL_AND2 A B Y vdd gnd
Xainv2 A A_n vdd gnd CMOS_INV
Xbinv2 B B_n vdd gnd CMOS_INV
Mpt_and and_int B A 0 0 CMOSN W={WN} L={2*LAMBDA}
Xbuf_and and_int Y vdd gnd CMOS_INV
.ends

* --- Domino CLA subckt (same as CMOS file) ---
.subckt DOMINO_C3_CLA G2 P2 G1 P1 G0 P0 C0 CLK Yout vdd gnd
M_footer eval CLK 0 0 CMOSN W={WN} L={2*LAMBDA}
M_pre dyn CLK vdd vdd CMOSP W={WP} L={2*LAMBDA}
M_keeper dyn Yout vdd vdd CMOSP W={WN} L={2*LAMBDA}

M_g2 dyn G2 eval eval CMOSN W={WN} L={2*LAMBDA}
M_p2g1_1 dyn P2 n1 eval CMOSN W={WN*2} L={2*LAMBDA}
M_p2g1_2 n1 G1 eval eval CMOSN W={WN*2} L={2*LAMBDA}
M_p2p1g0_1 dyn P2 n2 eval CMOSN W={WN*3} L={2*LAMBDA}
M_p2p1g0_2 n2 P1 n3 CMOSN W={WN*3} L={2*LAMBDA}
M_p2p1g0_3 n3 G0 eval eval CMOSN W={WN*3} L={2*LAMBDA}
M_p2p1p0c0_1 dyn P2 n4 eval CMOSN W={WN*4} L={2*LAMBDA}
M_p2p1p0c0_2 n4 P1 n5 CMOSN W={WN*4} L={2*LAMBDA}
M_p2p1p0c0_3 n5 P0 n6 CMOSN W={WN*4} L={2*LAMBDA}
M_p2p1p0c0_4 n6 C0 eval eval CMOSN W={WN*4} L={2*LAMBDA}

Xout_buf dyn Yout vdd gnd CMOS_INV
.ic V(dyn)= 'SUPPLY'
.ic V(n1)=0 V(n2)=0 V(n3)=0 V(n4)=0 V(n5)=0 V(n6)=0 V(eval)=0
.ends

* --- Instantiate CPL P/G blocks (true outputs used by domino) ---
Xp2 a2 b2 p2 vdd 0 CPL_XOR2
Xg2 a2 b2 g2 vdd 0 CPL_AND2
Xp1 a1 b1 p1 vdd 0 CPL_XOR2
Xg1 a1 b1 g1 vdd 0 CPL_AND2
Xp0 a0 b0 p0 vdd 0 CPL_XOR2
Xg0 a0 b0 g0 vdd 0 CPL_AND2

* Domino CLA instance (same)
Xc3 g2 p2 g1 p1 g0 p0 c0 clk c3_out vdd 0 DOMINO_C3_CLA

* load
Cload c3_out 0 10f

* --- Measurements ---
.meas tran t_rise TRIG v(c3_out) VAL='0.1*SUPPLY' RISE=1 TARG v(c3_out) VAL='0.9*SUPPLY' RISE=1
.meas tran t_fall TRIG v(c3_out) VAL='0.9*SUPPLY' FALL=1 TARG v(c3_out) VAL='0.1*SUPPLY' FALL=1
.meas tran energy PARAM='SUPPLY*ABS(INTEG(I(Vdd) from=0 to=160e-9))'
.meas tran avg_power PARAM='energy/160e-9'
.meas tran Ipeak MAX I(Vdd)

.control
set hcopypscolor=1
tran 0.1n 160n uic
run
plot v(clk) v(a2) v(b2) v(p2) v(g2) v(c3_out)
echo "t_rise = " $meas(t_rise)
echo "t_fall = " $meas(t_fall)
echo "energy = " $meas(energy)
echo "avg_power = " $meas(avg_power)
echo "Ipeak = " $meas(Ipeak)
.endc

.end
