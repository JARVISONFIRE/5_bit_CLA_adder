magic
tech scmos
timestamp 1764776976
<< nwell >>
rect 296 863 323 888
rect 242 809 267 832
rect 296 753 323 778
rect 252 661 277 684
rect 294 658 323 678
rect 294 653 321 658
rect 296 543 323 568
rect 296 432 323 457
rect 242 378 267 401
rect 296 322 323 347
rect 252 230 277 253
rect 294 227 323 247
rect 294 222 321 227
rect 296 112 323 137
rect 675 70 700 93
rect 710 69 742 89
rect 852 47 892 67
rect 905 47 930 70
rect 3 20 35 40
rect 46 20 70 40
rect 84 20 108 40
rect 122 21 147 44
rect 296 1 323 26
rect 675 -5 700 18
rect 710 -6 742 14
rect 3 -40 35 -20
rect 46 -40 70 -20
rect 84 -40 108 -20
rect 122 -39 147 -16
rect 242 -53 267 -30
rect 852 -31 892 -11
rect 905 -31 930 -8
rect 450 -64 482 -44
rect 492 -63 517 -43
rect 3 -100 35 -80
rect 46 -100 70 -80
rect 84 -100 108 -80
rect 122 -99 147 -76
rect 675 -80 700 -57
rect 710 -81 742 -61
rect 296 -109 323 -84
rect 455 -123 480 -100
rect 490 -124 522 -104
rect 852 -109 892 -89
rect 905 -109 930 -86
rect 3 -160 35 -140
rect 46 -160 70 -140
rect 84 -160 108 -140
rect 122 -159 147 -136
rect 675 -155 700 -132
rect 710 -156 742 -136
rect 3 -220 35 -200
rect 46 -220 70 -200
rect 84 -220 108 -200
rect 122 -219 147 -196
rect 252 -201 277 -178
rect 455 -183 480 -160
rect 490 -184 522 -164
rect 294 -204 323 -184
rect 852 -187 892 -167
rect 905 -187 930 -164
rect 294 -209 321 -204
rect 455 -243 480 -220
rect 490 -244 522 -224
rect 852 -265 892 -245
rect 905 -265 930 -242
rect 3 -290 35 -270
rect 46 -290 70 -270
rect 84 -290 108 -270
rect 122 -289 147 -266
rect 296 -319 323 -294
rect 455 -303 480 -280
rect 490 -304 522 -284
rect 3 -350 35 -330
rect 46 -350 70 -330
rect 84 -350 108 -330
rect 122 -349 147 -326
rect 3 -410 35 -390
rect 46 -410 70 -390
rect 84 -410 108 -390
rect 122 -409 147 -386
rect 296 -430 323 -405
rect 3 -470 35 -450
rect 46 -470 70 -450
rect 84 -470 108 -450
rect 122 -469 147 -446
rect 242 -484 267 -461
rect 3 -530 35 -510
rect 46 -530 70 -510
rect 84 -530 108 -510
rect 122 -529 147 -506
rect 296 -540 323 -515
rect 252 -632 277 -609
rect 294 -635 323 -615
rect 294 -640 321 -635
rect 296 -750 323 -725
rect 296 -861 323 -836
rect 242 -915 267 -892
rect 296 -971 323 -946
rect 252 -1063 277 -1040
rect 294 -1066 323 -1046
rect 294 -1071 321 -1066
rect 296 -1181 323 -1156
<< ntransistor >>
rect 308 842 310 850
rect 254 797 256 801
rect 308 732 310 740
rect 264 649 266 653
rect 308 632 310 640
rect 308 522 310 530
rect 308 411 310 419
rect 254 366 256 370
rect 308 301 310 309
rect 264 218 266 222
rect 308 201 310 209
rect 308 91 310 99
rect 686 58 688 62
rect 721 58 723 62
rect 729 58 731 62
rect 863 36 865 40
rect 871 36 873 40
rect 879 36 881 40
rect 917 35 919 39
rect 14 9 16 13
rect 57 9 59 13
rect 65 9 67 13
rect 95 9 97 13
rect 103 9 105 13
rect 134 9 136 13
rect 308 -20 310 -12
rect 686 -17 688 -13
rect 721 -17 723 -13
rect 729 -17 731 -13
rect 863 -42 865 -38
rect 871 -42 873 -38
rect 879 -42 881 -38
rect 14 -51 16 -47
rect 57 -51 59 -47
rect 65 -51 67 -47
rect 95 -51 97 -47
rect 103 -51 105 -47
rect 134 -51 136 -47
rect 917 -43 919 -39
rect 254 -65 256 -61
rect 461 -75 463 -71
rect 469 -75 471 -71
rect 504 -75 506 -71
rect 686 -92 688 -88
rect 721 -92 723 -88
rect 729 -92 731 -88
rect 14 -111 16 -107
rect 57 -111 59 -107
rect 65 -111 67 -107
rect 95 -111 97 -107
rect 103 -111 105 -107
rect 134 -111 136 -107
rect 308 -130 310 -122
rect 863 -120 865 -116
rect 871 -120 873 -116
rect 879 -120 881 -116
rect 466 -135 468 -131
rect 501 -135 503 -131
rect 509 -135 511 -131
rect 917 -121 919 -117
rect 14 -171 16 -167
rect 57 -171 59 -167
rect 65 -171 67 -167
rect 95 -171 97 -167
rect 103 -171 105 -167
rect 134 -171 136 -167
rect 686 -167 688 -163
rect 721 -167 723 -163
rect 729 -167 731 -163
rect 466 -195 468 -191
rect 501 -195 503 -191
rect 509 -195 511 -191
rect 863 -198 865 -194
rect 871 -198 873 -194
rect 879 -198 881 -194
rect 264 -213 266 -209
rect 917 -199 919 -195
rect 14 -231 16 -227
rect 57 -231 59 -227
rect 65 -231 67 -227
rect 95 -231 97 -227
rect 103 -231 105 -227
rect 134 -231 136 -227
rect 308 -230 310 -222
rect 466 -255 468 -251
rect 501 -255 503 -251
rect 509 -255 511 -251
rect 863 -276 865 -272
rect 871 -276 873 -272
rect 879 -276 881 -272
rect 14 -301 16 -297
rect 57 -301 59 -297
rect 65 -301 67 -297
rect 95 -301 97 -297
rect 103 -301 105 -297
rect 134 -301 136 -297
rect 917 -277 919 -273
rect 466 -315 468 -311
rect 501 -315 503 -311
rect 509 -315 511 -311
rect 308 -340 310 -332
rect 14 -361 16 -357
rect 57 -361 59 -357
rect 65 -361 67 -357
rect 95 -361 97 -357
rect 103 -361 105 -357
rect 134 -361 136 -357
rect 14 -421 16 -417
rect 57 -421 59 -417
rect 65 -421 67 -417
rect 95 -421 97 -417
rect 103 -421 105 -417
rect 134 -421 136 -417
rect 308 -451 310 -443
rect 14 -481 16 -477
rect 57 -481 59 -477
rect 65 -481 67 -477
rect 95 -481 97 -477
rect 103 -481 105 -477
rect 134 -481 136 -477
rect 254 -496 256 -492
rect 14 -541 16 -537
rect 57 -541 59 -537
rect 65 -541 67 -537
rect 95 -541 97 -537
rect 103 -541 105 -537
rect 134 -541 136 -537
rect 308 -561 310 -553
rect 264 -644 266 -640
rect 308 -661 310 -653
rect 308 -771 310 -763
rect 308 -882 310 -874
rect 254 -927 256 -923
rect 308 -992 310 -984
rect 264 -1075 266 -1071
rect 308 -1092 310 -1084
rect 308 -1202 310 -1194
<< ptransistor >>
rect 308 874 310 882
rect 254 816 256 824
rect 308 764 310 772
rect 264 668 266 676
rect 308 664 310 672
rect 308 554 310 562
rect 308 443 310 451
rect 254 385 256 393
rect 308 333 310 341
rect 264 237 266 245
rect 308 233 310 241
rect 308 123 310 131
rect 686 77 688 85
rect 721 75 723 83
rect 729 75 731 83
rect 863 53 865 61
rect 871 53 873 61
rect 879 53 881 61
rect 917 54 919 62
rect 14 26 16 34
rect 22 26 24 34
rect 57 26 59 34
rect 95 26 97 34
rect 134 28 136 36
rect 308 12 310 20
rect 686 2 688 10
rect 721 0 723 8
rect 729 0 731 8
rect 14 -34 16 -26
rect 22 -34 24 -26
rect 57 -34 59 -26
rect 95 -34 97 -26
rect 134 -32 136 -24
rect 863 -25 865 -17
rect 871 -25 873 -17
rect 879 -25 881 -17
rect 917 -24 919 -16
rect 254 -46 256 -38
rect 461 -58 463 -50
rect 469 -58 471 -50
rect 504 -56 506 -50
rect 686 -73 688 -65
rect 14 -94 16 -86
rect 22 -94 24 -86
rect 57 -94 59 -86
rect 95 -94 97 -86
rect 134 -92 136 -84
rect 721 -75 723 -67
rect 729 -75 731 -67
rect 308 -98 310 -90
rect 863 -103 865 -95
rect 871 -103 873 -95
rect 879 -103 881 -95
rect 917 -102 919 -94
rect 466 -116 468 -108
rect 501 -118 503 -110
rect 509 -118 511 -110
rect 14 -154 16 -146
rect 22 -154 24 -146
rect 57 -154 59 -146
rect 95 -154 97 -146
rect 134 -152 136 -144
rect 686 -148 688 -140
rect 721 -150 723 -142
rect 729 -150 731 -142
rect 466 -176 468 -168
rect 264 -194 266 -186
rect 14 -214 16 -206
rect 22 -214 24 -206
rect 57 -214 59 -206
rect 95 -214 97 -206
rect 134 -212 136 -204
rect 308 -198 310 -190
rect 501 -178 503 -170
rect 509 -178 511 -170
rect 863 -181 865 -173
rect 871 -181 873 -173
rect 879 -181 881 -173
rect 917 -180 919 -172
rect 466 -236 468 -228
rect 501 -238 503 -230
rect 509 -238 511 -230
rect 863 -259 865 -251
rect 871 -259 873 -251
rect 879 -259 881 -251
rect 917 -258 919 -250
rect 14 -284 16 -276
rect 22 -284 24 -276
rect 57 -284 59 -276
rect 95 -284 97 -276
rect 134 -282 136 -274
rect 466 -296 468 -288
rect 308 -308 310 -300
rect 501 -298 503 -290
rect 509 -298 511 -290
rect 14 -344 16 -336
rect 22 -344 24 -336
rect 57 -344 59 -336
rect 95 -344 97 -336
rect 134 -342 136 -334
rect 14 -404 16 -396
rect 22 -404 24 -396
rect 57 -404 59 -396
rect 95 -404 97 -396
rect 134 -402 136 -394
rect 308 -419 310 -411
rect 14 -464 16 -456
rect 22 -464 24 -456
rect 57 -464 59 -456
rect 95 -464 97 -456
rect 134 -462 136 -454
rect 254 -477 256 -469
rect 14 -524 16 -516
rect 22 -524 24 -516
rect 57 -524 59 -516
rect 95 -524 97 -516
rect 134 -522 136 -514
rect 308 -529 310 -521
rect 264 -625 266 -617
rect 308 -629 310 -621
rect 308 -739 310 -731
rect 308 -850 310 -842
rect 254 -908 256 -900
rect 308 -960 310 -952
rect 264 -1056 266 -1048
rect 308 -1060 310 -1052
rect 308 -1170 310 -1162
<< ndiffusion >>
rect 307 842 308 850
rect 310 842 311 850
rect 253 797 254 801
rect 256 797 257 801
rect 307 732 308 740
rect 310 732 311 740
rect 263 649 264 653
rect 266 649 267 653
rect 307 632 308 640
rect 310 632 311 640
rect 307 522 308 530
rect 310 522 311 530
rect 307 411 308 419
rect 310 411 311 419
rect 253 366 254 370
rect 256 366 257 370
rect 307 301 308 309
rect 310 301 311 309
rect 263 218 264 222
rect 266 218 267 222
rect 307 201 308 209
rect 310 201 311 209
rect 307 91 308 99
rect 310 91 311 99
rect 685 58 686 62
rect 688 58 689 62
rect 720 58 721 62
rect 723 58 724 62
rect 728 58 729 62
rect 731 58 732 62
rect 862 36 863 40
rect 865 36 866 40
rect 870 36 871 40
rect 873 36 874 40
rect 878 36 879 40
rect 881 36 882 40
rect 916 35 917 39
rect 919 35 920 39
rect 13 9 14 13
rect 16 9 17 13
rect 56 9 57 13
rect 59 9 60 13
rect 64 9 65 13
rect 67 9 68 13
rect 94 9 95 13
rect 97 9 98 13
rect 102 9 103 13
rect 105 9 106 13
rect 133 9 134 13
rect 136 9 137 13
rect 307 -20 308 -12
rect 310 -20 311 -12
rect 685 -17 686 -13
rect 688 -17 689 -13
rect 720 -17 721 -13
rect 723 -17 724 -13
rect 728 -17 729 -13
rect 731 -17 732 -13
rect 862 -42 863 -38
rect 865 -42 866 -38
rect 870 -42 871 -38
rect 873 -42 874 -38
rect 878 -42 879 -38
rect 881 -42 882 -38
rect 13 -51 14 -47
rect 16 -51 17 -47
rect 56 -51 57 -47
rect 59 -51 60 -47
rect 64 -51 65 -47
rect 67 -51 68 -47
rect 94 -51 95 -47
rect 97 -51 98 -47
rect 102 -51 103 -47
rect 105 -51 106 -47
rect 133 -51 134 -47
rect 136 -51 137 -47
rect 916 -43 917 -39
rect 919 -43 920 -39
rect 253 -65 254 -61
rect 256 -65 257 -61
rect 460 -75 461 -71
rect 463 -75 464 -71
rect 468 -75 469 -71
rect 471 -75 472 -71
rect 503 -75 504 -71
rect 506 -75 507 -71
rect 685 -92 686 -88
rect 688 -92 689 -88
rect 720 -92 721 -88
rect 723 -92 724 -88
rect 728 -92 729 -88
rect 731 -92 732 -88
rect 13 -111 14 -107
rect 16 -111 17 -107
rect 56 -111 57 -107
rect 59 -111 60 -107
rect 64 -111 65 -107
rect 67 -111 68 -107
rect 94 -111 95 -107
rect 97 -111 98 -107
rect 102 -111 103 -107
rect 105 -111 106 -107
rect 133 -111 134 -107
rect 136 -111 137 -107
rect 307 -130 308 -122
rect 310 -130 311 -122
rect 862 -120 863 -116
rect 865 -120 866 -116
rect 870 -120 871 -116
rect 873 -120 874 -116
rect 878 -120 879 -116
rect 881 -120 882 -116
rect 465 -135 466 -131
rect 468 -135 469 -131
rect 500 -135 501 -131
rect 503 -135 504 -131
rect 508 -135 509 -131
rect 511 -135 512 -131
rect 916 -121 917 -117
rect 919 -121 920 -117
rect 13 -171 14 -167
rect 16 -171 17 -167
rect 56 -171 57 -167
rect 59 -171 60 -167
rect 64 -171 65 -167
rect 67 -171 68 -167
rect 94 -171 95 -167
rect 97 -171 98 -167
rect 102 -171 103 -167
rect 105 -171 106 -167
rect 133 -171 134 -167
rect 136 -171 137 -167
rect 685 -167 686 -163
rect 688 -167 689 -163
rect 720 -167 721 -163
rect 723 -167 724 -163
rect 728 -167 729 -163
rect 731 -167 732 -163
rect 465 -195 466 -191
rect 468 -195 469 -191
rect 500 -195 501 -191
rect 503 -195 504 -191
rect 508 -195 509 -191
rect 511 -195 512 -191
rect 862 -198 863 -194
rect 865 -198 866 -194
rect 870 -198 871 -194
rect 873 -198 874 -194
rect 878 -198 879 -194
rect 881 -198 882 -194
rect 263 -213 264 -209
rect 266 -213 267 -209
rect 916 -199 917 -195
rect 919 -199 920 -195
rect 13 -231 14 -227
rect 16 -231 17 -227
rect 56 -231 57 -227
rect 59 -231 60 -227
rect 64 -231 65 -227
rect 67 -231 68 -227
rect 94 -231 95 -227
rect 97 -231 98 -227
rect 102 -231 103 -227
rect 105 -231 106 -227
rect 133 -231 134 -227
rect 136 -231 137 -227
rect 307 -230 308 -222
rect 310 -230 311 -222
rect 465 -255 466 -251
rect 468 -255 469 -251
rect 500 -255 501 -251
rect 503 -255 504 -251
rect 508 -255 509 -251
rect 511 -255 512 -251
rect 862 -276 863 -272
rect 865 -276 866 -272
rect 870 -276 871 -272
rect 873 -276 874 -272
rect 878 -276 879 -272
rect 881 -276 882 -272
rect 13 -301 14 -297
rect 16 -301 17 -297
rect 56 -301 57 -297
rect 59 -301 60 -297
rect 64 -301 65 -297
rect 67 -301 68 -297
rect 94 -301 95 -297
rect 97 -301 98 -297
rect 102 -301 103 -297
rect 105 -301 106 -297
rect 133 -301 134 -297
rect 136 -301 137 -297
rect 916 -277 917 -273
rect 919 -277 920 -273
rect 465 -315 466 -311
rect 468 -315 469 -311
rect 500 -315 501 -311
rect 503 -315 504 -311
rect 508 -315 509 -311
rect 511 -315 512 -311
rect 307 -340 308 -332
rect 310 -340 311 -332
rect 13 -361 14 -357
rect 16 -361 17 -357
rect 56 -361 57 -357
rect 59 -361 60 -357
rect 64 -361 65 -357
rect 67 -361 68 -357
rect 94 -361 95 -357
rect 97 -361 98 -357
rect 102 -361 103 -357
rect 105 -361 106 -357
rect 133 -361 134 -357
rect 136 -361 137 -357
rect 13 -421 14 -417
rect 16 -421 17 -417
rect 56 -421 57 -417
rect 59 -421 60 -417
rect 64 -421 65 -417
rect 67 -421 68 -417
rect 94 -421 95 -417
rect 97 -421 98 -417
rect 102 -421 103 -417
rect 105 -421 106 -417
rect 133 -421 134 -417
rect 136 -421 137 -417
rect 307 -451 308 -443
rect 310 -451 311 -443
rect 13 -481 14 -477
rect 16 -481 17 -477
rect 56 -481 57 -477
rect 59 -481 60 -477
rect 64 -481 65 -477
rect 67 -481 68 -477
rect 94 -481 95 -477
rect 97 -481 98 -477
rect 102 -481 103 -477
rect 105 -481 106 -477
rect 133 -481 134 -477
rect 136 -481 137 -477
rect 253 -496 254 -492
rect 256 -496 257 -492
rect 13 -541 14 -537
rect 16 -541 17 -537
rect 56 -541 57 -537
rect 59 -541 60 -537
rect 64 -541 65 -537
rect 67 -541 68 -537
rect 94 -541 95 -537
rect 97 -541 98 -537
rect 102 -541 103 -537
rect 105 -541 106 -537
rect 133 -541 134 -537
rect 136 -541 137 -537
rect 307 -561 308 -553
rect 310 -561 311 -553
rect 263 -644 264 -640
rect 266 -644 267 -640
rect 307 -661 308 -653
rect 310 -661 311 -653
rect 307 -771 308 -763
rect 310 -771 311 -763
rect 307 -882 308 -874
rect 310 -882 311 -874
rect 253 -927 254 -923
rect 256 -927 257 -923
rect 307 -992 308 -984
rect 310 -992 311 -984
rect 263 -1075 264 -1071
rect 266 -1075 267 -1071
rect 307 -1092 308 -1084
rect 310 -1092 311 -1084
rect 307 -1202 308 -1194
rect 310 -1202 311 -1194
<< pdiffusion >>
rect 307 874 308 882
rect 310 874 311 882
rect 253 816 254 824
rect 256 816 257 824
rect 307 764 308 772
rect 310 764 311 772
rect 263 668 264 676
rect 266 668 267 676
rect 307 664 308 672
rect 310 664 311 672
rect 307 554 308 562
rect 310 554 311 562
rect 307 443 308 451
rect 310 443 311 451
rect 253 385 254 393
rect 256 385 257 393
rect 307 333 308 341
rect 310 333 311 341
rect 263 237 264 245
rect 266 237 267 245
rect 307 233 308 241
rect 310 233 311 241
rect 307 123 308 131
rect 310 123 311 131
rect 685 77 686 85
rect 688 77 689 85
rect 720 75 721 83
rect 723 75 724 83
rect 728 75 729 83
rect 731 75 732 83
rect 862 53 863 61
rect 865 53 866 61
rect 870 53 871 61
rect 873 53 874 61
rect 878 53 879 61
rect 881 53 882 61
rect 916 54 917 62
rect 919 54 920 62
rect 13 26 14 34
rect 16 26 17 34
rect 21 26 22 34
rect 24 26 25 34
rect 56 26 57 34
rect 59 26 60 34
rect 94 26 95 34
rect 97 26 98 34
rect 133 28 134 36
rect 136 28 137 36
rect 307 12 308 20
rect 310 12 311 20
rect 685 2 686 10
rect 688 2 689 10
rect 720 0 721 8
rect 723 0 724 8
rect 728 0 729 8
rect 731 0 732 8
rect 13 -34 14 -26
rect 16 -34 17 -26
rect 21 -34 22 -26
rect 24 -34 25 -26
rect 56 -34 57 -26
rect 59 -34 60 -26
rect 94 -34 95 -26
rect 97 -34 98 -26
rect 133 -32 134 -24
rect 136 -32 137 -24
rect 862 -25 863 -17
rect 865 -25 866 -17
rect 870 -25 871 -17
rect 873 -25 874 -17
rect 878 -25 879 -17
rect 881 -25 882 -17
rect 916 -24 917 -16
rect 919 -24 920 -16
rect 253 -46 254 -38
rect 256 -46 257 -38
rect 460 -58 461 -50
rect 463 -58 464 -50
rect 468 -58 469 -50
rect 471 -58 472 -50
rect 503 -56 504 -50
rect 506 -56 507 -50
rect 685 -73 686 -65
rect 688 -73 689 -65
rect 13 -94 14 -86
rect 16 -94 17 -86
rect 21 -94 22 -86
rect 24 -94 25 -86
rect 56 -94 57 -86
rect 59 -94 60 -86
rect 94 -94 95 -86
rect 97 -94 98 -86
rect 133 -92 134 -84
rect 136 -92 137 -84
rect 720 -75 721 -67
rect 723 -75 724 -67
rect 728 -75 729 -67
rect 731 -75 732 -67
rect 307 -98 308 -90
rect 310 -98 311 -90
rect 862 -103 863 -95
rect 865 -103 866 -95
rect 870 -103 871 -95
rect 873 -103 874 -95
rect 878 -103 879 -95
rect 881 -103 882 -95
rect 916 -102 917 -94
rect 919 -102 920 -94
rect 465 -116 466 -108
rect 468 -116 469 -108
rect 500 -118 501 -110
rect 503 -118 504 -110
rect 508 -118 509 -110
rect 511 -118 512 -110
rect 13 -154 14 -146
rect 16 -154 17 -146
rect 21 -154 22 -146
rect 24 -154 25 -146
rect 56 -154 57 -146
rect 59 -154 60 -146
rect 94 -154 95 -146
rect 97 -154 98 -146
rect 133 -152 134 -144
rect 136 -152 137 -144
rect 685 -148 686 -140
rect 688 -148 689 -140
rect 720 -150 721 -142
rect 723 -150 724 -142
rect 728 -150 729 -142
rect 731 -150 732 -142
rect 465 -176 466 -168
rect 468 -176 469 -168
rect 263 -194 264 -186
rect 266 -194 267 -186
rect 13 -214 14 -206
rect 16 -214 17 -206
rect 21 -214 22 -206
rect 24 -214 25 -206
rect 56 -214 57 -206
rect 59 -214 60 -206
rect 94 -214 95 -206
rect 97 -214 98 -206
rect 133 -212 134 -204
rect 136 -212 137 -204
rect 307 -198 308 -190
rect 310 -198 311 -190
rect 500 -178 501 -170
rect 503 -178 504 -170
rect 508 -178 509 -170
rect 511 -178 512 -170
rect 862 -181 863 -173
rect 865 -181 866 -173
rect 870 -181 871 -173
rect 873 -181 874 -173
rect 878 -181 879 -173
rect 881 -181 882 -173
rect 916 -180 917 -172
rect 919 -180 920 -172
rect 465 -236 466 -228
rect 468 -236 469 -228
rect 500 -238 501 -230
rect 503 -238 504 -230
rect 508 -238 509 -230
rect 511 -238 512 -230
rect 862 -259 863 -251
rect 865 -259 866 -251
rect 870 -259 871 -251
rect 873 -259 874 -251
rect 878 -259 879 -251
rect 881 -259 882 -251
rect 916 -258 917 -250
rect 919 -258 920 -250
rect 13 -284 14 -276
rect 16 -284 17 -276
rect 21 -284 22 -276
rect 24 -284 25 -276
rect 56 -284 57 -276
rect 59 -284 60 -276
rect 94 -284 95 -276
rect 97 -284 98 -276
rect 133 -282 134 -274
rect 136 -282 137 -274
rect 465 -296 466 -288
rect 468 -296 469 -288
rect 307 -308 308 -300
rect 310 -308 311 -300
rect 500 -298 501 -290
rect 503 -298 504 -290
rect 508 -298 509 -290
rect 511 -298 512 -290
rect 13 -344 14 -336
rect 16 -344 17 -336
rect 21 -344 22 -336
rect 24 -344 25 -336
rect 56 -344 57 -336
rect 59 -344 60 -336
rect 94 -344 95 -336
rect 97 -344 98 -336
rect 133 -342 134 -334
rect 136 -342 137 -334
rect 13 -404 14 -396
rect 16 -404 17 -396
rect 21 -404 22 -396
rect 24 -404 25 -396
rect 56 -404 57 -396
rect 59 -404 60 -396
rect 94 -404 95 -396
rect 97 -404 98 -396
rect 133 -402 134 -394
rect 136 -402 137 -394
rect 307 -419 308 -411
rect 310 -419 311 -411
rect 13 -464 14 -456
rect 16 -464 17 -456
rect 21 -464 22 -456
rect 24 -464 25 -456
rect 56 -464 57 -456
rect 59 -464 60 -456
rect 94 -464 95 -456
rect 97 -464 98 -456
rect 133 -462 134 -454
rect 136 -462 137 -454
rect 253 -477 254 -469
rect 256 -477 257 -469
rect 13 -524 14 -516
rect 16 -524 17 -516
rect 21 -524 22 -516
rect 24 -524 25 -516
rect 56 -524 57 -516
rect 59 -524 60 -516
rect 94 -524 95 -516
rect 97 -524 98 -516
rect 133 -522 134 -514
rect 136 -522 137 -514
rect 307 -529 308 -521
rect 310 -529 311 -521
rect 263 -625 264 -617
rect 266 -625 267 -617
rect 307 -629 308 -621
rect 310 -629 311 -621
rect 307 -739 308 -731
rect 310 -739 311 -731
rect 307 -850 308 -842
rect 310 -850 311 -842
rect 253 -908 254 -900
rect 256 -908 257 -900
rect 307 -960 308 -952
rect 310 -960 311 -952
rect 263 -1056 264 -1048
rect 266 -1056 267 -1048
rect 307 -1060 308 -1052
rect 310 -1060 311 -1052
rect 307 -1170 308 -1162
rect 310 -1170 311 -1162
<< ndcontact >>
rect 303 842 307 850
rect 311 842 315 850
rect 249 797 253 801
rect 257 797 261 801
rect 303 732 307 740
rect 311 732 315 740
rect 259 649 263 653
rect 267 649 271 653
rect 303 632 307 640
rect 311 632 315 640
rect 303 522 307 530
rect 311 522 315 530
rect 303 411 307 419
rect 311 411 315 419
rect 249 366 253 370
rect 257 366 261 370
rect 303 301 307 309
rect 311 301 315 309
rect 259 218 263 222
rect 267 218 271 222
rect 303 201 307 209
rect 311 201 315 209
rect 303 91 307 99
rect 311 91 315 99
rect 681 58 685 62
rect 689 58 693 62
rect 716 58 720 62
rect 724 58 728 62
rect 732 58 736 62
rect 858 36 862 40
rect 866 36 870 40
rect 874 36 878 40
rect 882 36 886 40
rect 912 35 916 39
rect 920 35 924 39
rect 9 9 13 13
rect 17 9 21 13
rect 52 9 56 13
rect 60 9 64 13
rect 68 9 72 13
rect 90 9 94 13
rect 98 9 102 13
rect 106 9 110 13
rect 129 9 133 13
rect 137 9 141 13
rect 303 -20 307 -12
rect 311 -20 315 -12
rect 681 -17 685 -13
rect 689 -17 693 -13
rect 716 -17 720 -13
rect 724 -17 728 -13
rect 732 -17 736 -13
rect 858 -42 862 -38
rect 866 -42 870 -38
rect 874 -42 878 -38
rect 882 -42 886 -38
rect 9 -51 13 -47
rect 17 -51 21 -47
rect 52 -51 56 -47
rect 60 -51 64 -47
rect 68 -51 72 -47
rect 90 -51 94 -47
rect 98 -51 102 -47
rect 106 -51 110 -47
rect 129 -51 133 -47
rect 137 -51 141 -47
rect 912 -43 916 -39
rect 920 -43 924 -39
rect 249 -65 253 -61
rect 257 -65 261 -61
rect 456 -75 460 -71
rect 464 -75 468 -71
rect 472 -75 476 -71
rect 499 -75 503 -71
rect 507 -75 511 -71
rect 681 -92 685 -88
rect 689 -92 693 -88
rect 716 -92 720 -88
rect 724 -92 728 -88
rect 732 -92 736 -88
rect 9 -111 13 -107
rect 17 -111 21 -107
rect 52 -111 56 -107
rect 60 -111 64 -107
rect 68 -111 72 -107
rect 90 -111 94 -107
rect 98 -111 102 -107
rect 106 -111 110 -107
rect 129 -111 133 -107
rect 137 -111 141 -107
rect 303 -130 307 -122
rect 311 -130 315 -122
rect 858 -120 862 -116
rect 866 -120 870 -116
rect 874 -120 878 -116
rect 882 -120 886 -116
rect 461 -135 465 -131
rect 469 -135 473 -131
rect 496 -135 500 -131
rect 504 -135 508 -131
rect 512 -135 516 -131
rect 912 -121 916 -117
rect 920 -121 924 -117
rect 9 -171 13 -167
rect 17 -171 21 -167
rect 52 -171 56 -167
rect 60 -171 64 -167
rect 68 -171 72 -167
rect 90 -171 94 -167
rect 98 -171 102 -167
rect 106 -171 110 -167
rect 129 -171 133 -167
rect 137 -171 141 -167
rect 681 -167 685 -163
rect 689 -167 693 -163
rect 716 -167 720 -163
rect 724 -167 728 -163
rect 732 -167 736 -163
rect 461 -195 465 -191
rect 469 -195 473 -191
rect 496 -195 500 -191
rect 504 -195 508 -191
rect 512 -195 516 -191
rect 858 -198 862 -194
rect 866 -198 870 -194
rect 874 -198 878 -194
rect 882 -198 886 -194
rect 259 -213 263 -209
rect 267 -213 271 -209
rect 912 -199 916 -195
rect 920 -199 924 -195
rect 9 -231 13 -227
rect 17 -231 21 -227
rect 52 -231 56 -227
rect 60 -231 64 -227
rect 68 -231 72 -227
rect 90 -231 94 -227
rect 98 -231 102 -227
rect 106 -231 110 -227
rect 129 -231 133 -227
rect 137 -231 141 -227
rect 303 -230 307 -222
rect 311 -230 315 -222
rect 461 -255 465 -251
rect 469 -255 473 -251
rect 496 -255 500 -251
rect 504 -255 508 -251
rect 512 -255 516 -251
rect 858 -276 862 -272
rect 866 -276 870 -272
rect 874 -276 878 -272
rect 882 -276 886 -272
rect 9 -301 13 -297
rect 17 -301 21 -297
rect 52 -301 56 -297
rect 60 -301 64 -297
rect 68 -301 72 -297
rect 90 -301 94 -297
rect 98 -301 102 -297
rect 106 -301 110 -297
rect 129 -301 133 -297
rect 137 -301 141 -297
rect 912 -277 916 -273
rect 920 -277 924 -273
rect 461 -315 465 -311
rect 469 -315 473 -311
rect 496 -315 500 -311
rect 504 -315 508 -311
rect 512 -315 516 -311
rect 303 -340 307 -332
rect 311 -340 315 -332
rect 9 -361 13 -357
rect 17 -361 21 -357
rect 52 -361 56 -357
rect 60 -361 64 -357
rect 68 -361 72 -357
rect 90 -361 94 -357
rect 98 -361 102 -357
rect 106 -361 110 -357
rect 129 -361 133 -357
rect 137 -361 141 -357
rect 9 -421 13 -417
rect 17 -421 21 -417
rect 52 -421 56 -417
rect 60 -421 64 -417
rect 68 -421 72 -417
rect 90 -421 94 -417
rect 98 -421 102 -417
rect 106 -421 110 -417
rect 129 -421 133 -417
rect 137 -421 141 -417
rect 303 -451 307 -443
rect 311 -451 315 -443
rect 9 -481 13 -477
rect 17 -481 21 -477
rect 52 -481 56 -477
rect 60 -481 64 -477
rect 68 -481 72 -477
rect 90 -481 94 -477
rect 98 -481 102 -477
rect 106 -481 110 -477
rect 129 -481 133 -477
rect 137 -481 141 -477
rect 249 -496 253 -492
rect 257 -496 261 -492
rect 9 -541 13 -537
rect 17 -541 21 -537
rect 52 -541 56 -537
rect 60 -541 64 -537
rect 68 -541 72 -537
rect 90 -541 94 -537
rect 98 -541 102 -537
rect 106 -541 110 -537
rect 129 -541 133 -537
rect 137 -541 141 -537
rect 303 -561 307 -553
rect 311 -561 315 -553
rect 259 -644 263 -640
rect 267 -644 271 -640
rect 303 -661 307 -653
rect 311 -661 315 -653
rect 303 -771 307 -763
rect 311 -771 315 -763
rect 303 -882 307 -874
rect 311 -882 315 -874
rect 249 -927 253 -923
rect 257 -927 261 -923
rect 303 -992 307 -984
rect 311 -992 315 -984
rect 259 -1075 263 -1071
rect 267 -1075 271 -1071
rect 303 -1092 307 -1084
rect 311 -1092 315 -1084
rect 303 -1202 307 -1194
rect 311 -1202 315 -1194
<< pdcontact >>
rect 303 874 307 882
rect 311 874 315 882
rect 249 816 253 824
rect 257 816 261 824
rect 303 764 307 772
rect 311 764 315 772
rect 259 668 263 676
rect 267 668 271 676
rect 303 664 307 672
rect 311 664 315 672
rect 303 554 307 562
rect 311 554 315 562
rect 303 443 307 451
rect 311 443 315 451
rect 249 385 253 393
rect 257 385 261 393
rect 303 333 307 341
rect 311 333 315 341
rect 259 237 263 245
rect 267 237 271 245
rect 303 233 307 241
rect 311 233 315 241
rect 303 123 307 131
rect 311 123 315 131
rect 681 77 685 85
rect 689 77 693 85
rect 716 75 720 83
rect 724 75 728 83
rect 732 75 736 83
rect 858 53 862 61
rect 866 53 870 61
rect 874 53 878 61
rect 882 53 886 61
rect 912 54 916 62
rect 920 54 924 62
rect 9 26 13 34
rect 17 26 21 34
rect 25 26 29 34
rect 52 26 56 34
rect 60 26 64 34
rect 90 26 94 34
rect 98 26 102 34
rect 129 28 133 36
rect 137 28 141 36
rect 303 12 307 20
rect 311 12 315 20
rect 681 2 685 10
rect 689 2 693 10
rect 716 0 720 8
rect 724 0 728 8
rect 732 0 736 8
rect 9 -34 13 -26
rect 17 -34 21 -26
rect 25 -34 29 -26
rect 52 -34 56 -26
rect 60 -34 64 -26
rect 90 -34 94 -26
rect 98 -34 102 -26
rect 129 -32 133 -24
rect 137 -32 141 -24
rect 858 -25 862 -17
rect 866 -25 870 -17
rect 874 -25 878 -17
rect 882 -25 886 -17
rect 912 -24 916 -16
rect 920 -24 924 -16
rect 249 -46 253 -38
rect 257 -46 261 -38
rect 456 -58 460 -50
rect 464 -58 468 -50
rect 472 -58 476 -50
rect 499 -56 503 -50
rect 507 -56 511 -50
rect 681 -73 685 -65
rect 689 -73 693 -65
rect 9 -94 13 -86
rect 17 -94 21 -86
rect 25 -94 29 -86
rect 52 -94 56 -86
rect 60 -94 64 -86
rect 90 -94 94 -86
rect 98 -94 102 -86
rect 129 -92 133 -84
rect 137 -92 141 -84
rect 716 -75 720 -67
rect 724 -75 728 -67
rect 732 -75 736 -67
rect 303 -98 307 -90
rect 311 -98 315 -90
rect 858 -103 862 -95
rect 866 -103 870 -95
rect 874 -103 878 -95
rect 882 -103 886 -95
rect 912 -102 916 -94
rect 920 -102 924 -94
rect 461 -116 465 -108
rect 469 -116 473 -108
rect 496 -118 500 -110
rect 504 -118 508 -110
rect 512 -118 516 -110
rect 9 -154 13 -146
rect 17 -154 21 -146
rect 25 -154 29 -146
rect 52 -154 56 -146
rect 60 -154 64 -146
rect 90 -154 94 -146
rect 98 -154 102 -146
rect 129 -152 133 -144
rect 137 -152 141 -144
rect 681 -148 685 -140
rect 689 -148 693 -140
rect 716 -150 720 -142
rect 724 -150 728 -142
rect 732 -150 736 -142
rect 461 -176 465 -168
rect 469 -176 473 -168
rect 259 -194 263 -186
rect 267 -194 271 -186
rect 9 -214 13 -206
rect 17 -214 21 -206
rect 25 -214 29 -206
rect 52 -214 56 -206
rect 60 -214 64 -206
rect 90 -214 94 -206
rect 98 -214 102 -206
rect 129 -212 133 -204
rect 137 -212 141 -204
rect 303 -198 307 -190
rect 311 -198 315 -190
rect 496 -178 500 -170
rect 504 -178 508 -170
rect 512 -178 516 -170
rect 858 -181 862 -173
rect 866 -181 870 -173
rect 874 -181 878 -173
rect 882 -181 886 -173
rect 912 -180 916 -172
rect 920 -180 924 -172
rect 461 -236 465 -228
rect 469 -236 473 -228
rect 496 -238 500 -230
rect 504 -238 508 -230
rect 512 -238 516 -230
rect 858 -259 862 -251
rect 866 -259 870 -251
rect 874 -259 878 -251
rect 882 -259 886 -251
rect 912 -258 916 -250
rect 920 -258 924 -250
rect 9 -284 13 -276
rect 17 -284 21 -276
rect 25 -284 29 -276
rect 52 -284 56 -276
rect 60 -284 64 -276
rect 90 -284 94 -276
rect 98 -284 102 -276
rect 129 -282 133 -274
rect 137 -282 141 -274
rect 461 -296 465 -288
rect 469 -296 473 -288
rect 303 -308 307 -300
rect 311 -308 315 -300
rect 496 -298 500 -290
rect 504 -298 508 -290
rect 512 -298 516 -290
rect 9 -344 13 -336
rect 17 -344 21 -336
rect 25 -344 29 -336
rect 52 -344 56 -336
rect 60 -344 64 -336
rect 90 -344 94 -336
rect 98 -344 102 -336
rect 129 -342 133 -334
rect 137 -342 141 -334
rect 9 -404 13 -396
rect 17 -404 21 -396
rect 25 -404 29 -396
rect 52 -404 56 -396
rect 60 -404 64 -396
rect 90 -404 94 -396
rect 98 -404 102 -396
rect 129 -402 133 -394
rect 137 -402 141 -394
rect 303 -419 307 -411
rect 311 -419 315 -411
rect 9 -464 13 -456
rect 17 -464 21 -456
rect 25 -464 29 -456
rect 52 -464 56 -456
rect 60 -464 64 -456
rect 90 -464 94 -456
rect 98 -464 102 -456
rect 129 -462 133 -454
rect 137 -462 141 -454
rect 249 -477 253 -469
rect 257 -477 261 -469
rect 9 -524 13 -516
rect 17 -524 21 -516
rect 25 -524 29 -516
rect 52 -524 56 -516
rect 60 -524 64 -516
rect 90 -524 94 -516
rect 98 -524 102 -516
rect 129 -522 133 -514
rect 137 -522 141 -514
rect 303 -529 307 -521
rect 311 -529 315 -521
rect 259 -625 263 -617
rect 267 -625 271 -617
rect 303 -629 307 -621
rect 311 -629 315 -621
rect 303 -739 307 -731
rect 311 -739 315 -731
rect 303 -850 307 -842
rect 311 -850 315 -842
rect 249 -908 253 -900
rect 257 -908 261 -900
rect 303 -960 307 -952
rect 311 -960 315 -952
rect 259 -1056 263 -1048
rect 267 -1056 271 -1048
rect 303 -1060 307 -1052
rect 311 -1060 315 -1052
rect 303 -1170 307 -1162
rect 311 -1170 315 -1162
<< nsubstratencontact >>
rect 315 866 319 870
rect 315 756 319 760
rect 314 656 318 660
rect 315 546 319 550
rect 315 435 319 439
rect 315 325 319 329
rect 314 225 318 229
rect 315 115 319 119
rect 315 4 319 8
rect 315 -106 319 -102
rect 314 -206 318 -202
rect 315 -316 319 -312
rect 315 -427 319 -423
rect 315 -537 319 -533
rect 314 -637 318 -633
rect 315 -747 319 -743
rect 315 -858 319 -854
rect 315 -968 319 -964
rect 314 -1068 318 -1064
rect 315 -1178 319 -1174
<< polysilicon >>
rect 308 882 310 889
rect 308 868 310 874
rect 308 850 310 856
rect 308 839 310 842
rect 254 824 256 827
rect 254 801 256 816
rect 254 794 256 797
rect 308 772 310 780
rect 308 758 310 764
rect 308 740 310 746
rect 308 728 310 732
rect 264 676 266 679
rect 308 672 310 679
rect 264 653 266 668
rect 308 658 310 664
rect 264 646 266 649
rect 308 640 310 646
rect 308 628 310 632
rect 308 562 310 569
rect 308 548 310 554
rect 308 530 310 536
rect 308 518 310 522
rect 308 451 310 458
rect 308 437 310 443
rect 308 419 310 425
rect 308 408 310 411
rect 254 393 256 396
rect 254 370 256 385
rect 254 363 256 366
rect 308 341 310 349
rect 308 327 310 333
rect 308 309 310 315
rect 308 297 310 301
rect 264 245 266 248
rect 308 241 310 248
rect 264 222 266 237
rect 308 227 310 233
rect 264 215 266 218
rect 308 209 310 215
rect 308 197 310 201
rect 308 131 310 138
rect 308 117 310 123
rect 308 99 310 105
rect 308 87 310 91
rect 686 85 688 88
rect 721 83 723 87
rect 729 83 731 87
rect 686 62 688 77
rect 721 65 723 75
rect 711 63 723 65
rect 711 62 713 63
rect 721 62 723 63
rect 729 62 731 75
rect 863 61 865 65
rect 871 61 873 65
rect 879 61 881 65
rect 917 62 919 65
rect 686 55 688 58
rect 721 54 723 58
rect 729 54 731 58
rect 863 43 865 53
rect 855 41 865 43
rect 863 40 865 41
rect 871 40 873 53
rect 879 49 881 53
rect 879 47 896 49
rect 879 40 881 47
rect 14 34 16 38
rect 22 36 32 38
rect 22 34 24 36
rect 57 34 59 38
rect 95 34 97 38
rect 134 36 136 39
rect 917 39 919 54
rect 863 32 865 36
rect 14 21 16 26
rect 22 23 24 26
rect 57 20 59 26
rect 95 20 97 26
rect 14 13 16 17
rect 57 13 59 16
rect 65 15 75 17
rect 65 13 67 15
rect 95 13 97 16
rect 103 15 113 17
rect 103 13 105 15
rect 134 13 136 28
rect 308 20 310 27
rect 871 24 873 36
rect 879 32 881 36
rect 917 32 919 35
rect 14 5 16 9
rect 57 5 59 9
rect 65 5 67 9
rect 95 5 97 9
rect 103 5 105 9
rect 134 6 136 9
rect 308 6 310 12
rect 686 10 688 13
rect 721 8 723 12
rect 729 8 731 12
rect 308 -12 310 -6
rect 686 -13 688 2
rect 721 -10 723 0
rect 711 -12 723 -10
rect 711 -13 713 -12
rect 721 -13 723 -12
rect 729 -13 731 0
rect 863 -17 865 -13
rect 871 -17 873 -13
rect 879 -17 881 -13
rect 917 -16 919 -13
rect 686 -20 688 -17
rect 14 -26 16 -22
rect 22 -24 32 -22
rect 22 -26 24 -24
rect 57 -26 59 -22
rect 95 -26 97 -22
rect 134 -24 136 -21
rect 308 -23 310 -20
rect 721 -21 723 -17
rect 729 -21 731 -17
rect 14 -39 16 -34
rect 22 -37 24 -34
rect 57 -40 59 -34
rect 95 -40 97 -34
rect 14 -47 16 -43
rect 57 -47 59 -44
rect 65 -45 75 -43
rect 65 -47 67 -45
rect 95 -47 97 -44
rect 103 -45 113 -43
rect 103 -47 105 -45
rect 134 -47 136 -32
rect 863 -35 865 -25
rect 254 -38 256 -35
rect 855 -37 865 -35
rect 863 -38 865 -37
rect 871 -38 873 -25
rect 879 -29 881 -25
rect 879 -31 896 -29
rect 879 -38 881 -31
rect 917 -39 919 -24
rect 14 -55 16 -51
rect 57 -55 59 -51
rect 65 -55 67 -51
rect 95 -55 97 -51
rect 103 -55 105 -51
rect 134 -54 136 -51
rect 254 -61 256 -46
rect 461 -50 463 -46
rect 469 -50 471 -46
rect 504 -50 506 -44
rect 863 -46 865 -42
rect 871 -54 873 -42
rect 879 -46 881 -42
rect 917 -46 919 -43
rect 254 -68 256 -65
rect 461 -71 463 -58
rect 469 -68 471 -58
rect 469 -70 481 -68
rect 469 -71 471 -70
rect 479 -71 481 -70
rect 504 -71 506 -56
rect 686 -65 688 -62
rect 721 -67 723 -63
rect 729 -67 731 -63
rect 14 -86 16 -82
rect 22 -84 32 -82
rect 22 -86 24 -84
rect 57 -86 59 -82
rect 95 -86 97 -82
rect 134 -84 136 -81
rect 461 -79 463 -75
rect 469 -79 471 -75
rect 504 -78 506 -75
rect 308 -90 310 -82
rect 686 -88 688 -73
rect 721 -85 723 -75
rect 711 -87 723 -85
rect 711 -88 713 -87
rect 721 -88 723 -87
rect 729 -88 731 -75
rect 14 -99 16 -94
rect 22 -97 24 -94
rect 57 -100 59 -94
rect 95 -100 97 -94
rect 14 -107 16 -103
rect 57 -107 59 -104
rect 65 -105 75 -103
rect 65 -107 67 -105
rect 95 -107 97 -104
rect 103 -105 113 -103
rect 103 -107 105 -105
rect 134 -107 136 -92
rect 686 -95 688 -92
rect 721 -96 723 -92
rect 729 -96 731 -92
rect 863 -95 865 -91
rect 871 -95 873 -91
rect 879 -95 881 -91
rect 917 -94 919 -91
rect 308 -104 310 -98
rect 466 -108 468 -105
rect 14 -115 16 -111
rect 57 -115 59 -111
rect 65 -115 67 -111
rect 95 -115 97 -111
rect 103 -115 105 -111
rect 134 -114 136 -111
rect 501 -110 503 -106
rect 509 -110 511 -106
rect 308 -122 310 -116
rect 308 -134 310 -130
rect 466 -131 468 -116
rect 863 -113 865 -103
rect 855 -115 865 -113
rect 863 -116 865 -115
rect 871 -116 873 -103
rect 879 -107 881 -103
rect 879 -109 896 -107
rect 879 -116 881 -109
rect 501 -128 503 -118
rect 491 -130 503 -128
rect 491 -131 493 -130
rect 501 -131 503 -130
rect 509 -131 511 -118
rect 917 -117 919 -102
rect 863 -124 865 -120
rect 871 -132 873 -120
rect 879 -124 881 -120
rect 917 -124 919 -121
rect 466 -138 468 -135
rect 501 -139 503 -135
rect 509 -139 511 -135
rect 686 -140 688 -137
rect 14 -146 16 -142
rect 22 -144 32 -142
rect 22 -146 24 -144
rect 57 -146 59 -142
rect 95 -146 97 -142
rect 134 -144 136 -141
rect 721 -142 723 -138
rect 729 -142 731 -138
rect 14 -159 16 -154
rect 22 -157 24 -154
rect 57 -160 59 -154
rect 95 -160 97 -154
rect 14 -167 16 -163
rect 57 -167 59 -164
rect 65 -165 75 -163
rect 65 -167 67 -165
rect 95 -167 97 -164
rect 103 -165 113 -163
rect 103 -167 105 -165
rect 134 -167 136 -152
rect 686 -163 688 -148
rect 721 -160 723 -150
rect 711 -162 723 -160
rect 711 -163 713 -162
rect 721 -163 723 -162
rect 729 -163 731 -150
rect 466 -168 468 -165
rect 14 -175 16 -171
rect 57 -175 59 -171
rect 65 -175 67 -171
rect 95 -175 97 -171
rect 103 -175 105 -171
rect 134 -174 136 -171
rect 501 -170 503 -166
rect 509 -170 511 -166
rect 686 -170 688 -167
rect 264 -186 266 -183
rect 308 -190 310 -183
rect 14 -206 16 -202
rect 22 -204 32 -202
rect 22 -206 24 -204
rect 57 -206 59 -202
rect 95 -206 97 -202
rect 134 -204 136 -201
rect 264 -209 266 -194
rect 466 -191 468 -176
rect 721 -171 723 -167
rect 729 -171 731 -167
rect 863 -173 865 -169
rect 871 -173 873 -169
rect 879 -173 881 -169
rect 917 -172 919 -169
rect 501 -188 503 -178
rect 491 -190 503 -188
rect 491 -191 493 -190
rect 501 -191 503 -190
rect 509 -191 511 -178
rect 863 -191 865 -181
rect 855 -193 865 -191
rect 863 -194 865 -193
rect 871 -194 873 -181
rect 879 -185 881 -181
rect 879 -187 896 -185
rect 879 -194 881 -187
rect 466 -198 468 -195
rect 308 -204 310 -198
rect 501 -199 503 -195
rect 509 -199 511 -195
rect 917 -195 919 -180
rect 863 -202 865 -198
rect 14 -219 16 -214
rect 22 -217 24 -214
rect 57 -220 59 -214
rect 95 -220 97 -214
rect 14 -227 16 -223
rect 57 -227 59 -224
rect 65 -225 75 -223
rect 65 -227 67 -225
rect 95 -227 97 -224
rect 103 -225 113 -223
rect 103 -227 105 -225
rect 134 -227 136 -212
rect 871 -210 873 -198
rect 879 -202 881 -198
rect 917 -202 919 -199
rect 264 -216 266 -213
rect 308 -222 310 -216
rect 466 -228 468 -225
rect 14 -235 16 -231
rect 57 -235 59 -231
rect 65 -235 67 -231
rect 95 -235 97 -231
rect 103 -235 105 -231
rect 134 -234 136 -231
rect 308 -234 310 -230
rect 501 -230 503 -226
rect 509 -230 511 -226
rect 466 -251 468 -236
rect 501 -248 503 -238
rect 491 -250 503 -248
rect 491 -251 493 -250
rect 501 -251 503 -250
rect 509 -251 511 -238
rect 863 -251 865 -247
rect 871 -251 873 -247
rect 879 -251 881 -247
rect 917 -250 919 -247
rect 466 -258 468 -255
rect 501 -259 503 -255
rect 509 -259 511 -255
rect 863 -269 865 -259
rect 14 -276 16 -272
rect 22 -274 32 -272
rect 22 -276 24 -274
rect 57 -276 59 -272
rect 95 -276 97 -272
rect 134 -274 136 -271
rect 855 -271 865 -269
rect 863 -272 865 -271
rect 871 -272 873 -259
rect 879 -263 881 -259
rect 879 -265 896 -263
rect 879 -272 881 -265
rect 917 -273 919 -258
rect 863 -280 865 -276
rect 14 -289 16 -284
rect 22 -287 24 -284
rect 57 -290 59 -284
rect 95 -290 97 -284
rect 14 -297 16 -293
rect 57 -297 59 -294
rect 65 -295 75 -293
rect 65 -297 67 -295
rect 95 -297 97 -294
rect 103 -295 113 -293
rect 103 -297 105 -295
rect 134 -297 136 -282
rect 466 -288 468 -285
rect 308 -300 310 -293
rect 501 -290 503 -286
rect 509 -290 511 -286
rect 871 -288 873 -276
rect 879 -280 881 -276
rect 917 -280 919 -277
rect 14 -305 16 -301
rect 57 -305 59 -301
rect 65 -305 67 -301
rect 95 -305 97 -301
rect 103 -305 105 -301
rect 134 -304 136 -301
rect 308 -314 310 -308
rect 466 -311 468 -296
rect 501 -308 503 -298
rect 491 -310 503 -308
rect 491 -311 493 -310
rect 501 -311 503 -310
rect 509 -311 511 -298
rect 466 -318 468 -315
rect 501 -319 503 -315
rect 509 -319 511 -315
rect 14 -336 16 -332
rect 22 -334 32 -332
rect 22 -336 24 -334
rect 57 -336 59 -332
rect 95 -336 97 -332
rect 134 -334 136 -331
rect 308 -332 310 -326
rect 14 -349 16 -344
rect 22 -347 24 -344
rect 57 -350 59 -344
rect 95 -350 97 -344
rect 14 -357 16 -353
rect 57 -357 59 -354
rect 65 -355 75 -353
rect 65 -357 67 -355
rect 95 -357 97 -354
rect 103 -355 113 -353
rect 103 -357 105 -355
rect 134 -357 136 -342
rect 308 -344 310 -340
rect 14 -365 16 -361
rect 57 -365 59 -361
rect 65 -365 67 -361
rect 95 -365 97 -361
rect 103 -365 105 -361
rect 134 -364 136 -361
rect 14 -396 16 -392
rect 22 -394 32 -392
rect 22 -396 24 -394
rect 57 -396 59 -392
rect 95 -396 97 -392
rect 134 -394 136 -391
rect 14 -409 16 -404
rect 22 -407 24 -404
rect 57 -410 59 -404
rect 95 -410 97 -404
rect 14 -417 16 -413
rect 57 -417 59 -414
rect 65 -415 75 -413
rect 65 -417 67 -415
rect 95 -417 97 -414
rect 103 -415 113 -413
rect 103 -417 105 -415
rect 134 -417 136 -402
rect 308 -411 310 -404
rect 14 -425 16 -421
rect 57 -425 59 -421
rect 65 -425 67 -421
rect 95 -425 97 -421
rect 103 -425 105 -421
rect 134 -424 136 -421
rect 308 -425 310 -419
rect 308 -443 310 -437
rect 14 -456 16 -452
rect 22 -454 32 -452
rect 22 -456 24 -454
rect 57 -456 59 -452
rect 95 -456 97 -452
rect 134 -454 136 -451
rect 308 -454 310 -451
rect 14 -469 16 -464
rect 22 -467 24 -464
rect 57 -470 59 -464
rect 95 -470 97 -464
rect 14 -477 16 -473
rect 57 -477 59 -474
rect 65 -475 75 -473
rect 65 -477 67 -475
rect 95 -477 97 -474
rect 103 -475 113 -473
rect 103 -477 105 -475
rect 134 -477 136 -462
rect 254 -469 256 -466
rect 14 -485 16 -481
rect 57 -485 59 -481
rect 65 -485 67 -481
rect 95 -485 97 -481
rect 103 -485 105 -481
rect 134 -484 136 -481
rect 254 -492 256 -477
rect 254 -499 256 -496
rect 14 -516 16 -512
rect 22 -514 32 -512
rect 22 -516 24 -514
rect 57 -516 59 -512
rect 95 -516 97 -512
rect 134 -514 136 -511
rect 308 -521 310 -513
rect 14 -529 16 -524
rect 22 -527 24 -524
rect 57 -530 59 -524
rect 95 -530 97 -524
rect 14 -537 16 -533
rect 57 -537 59 -534
rect 65 -535 75 -533
rect 65 -537 67 -535
rect 95 -537 97 -534
rect 103 -535 113 -533
rect 103 -537 105 -535
rect 134 -537 136 -522
rect 308 -535 310 -529
rect 14 -545 16 -541
rect 57 -545 59 -541
rect 65 -545 67 -541
rect 95 -545 97 -541
rect 103 -545 105 -541
rect 134 -544 136 -541
rect 308 -553 310 -547
rect 308 -565 310 -561
rect 264 -617 266 -614
rect 308 -621 310 -614
rect 264 -640 266 -625
rect 308 -635 310 -629
rect 264 -647 266 -644
rect 308 -653 310 -647
rect 308 -665 310 -661
rect 308 -731 310 -724
rect 308 -745 310 -739
rect 308 -763 310 -757
rect 308 -775 310 -771
rect 308 -842 310 -835
rect 308 -856 310 -850
rect 308 -874 310 -868
rect 308 -885 310 -882
rect 254 -900 256 -897
rect 254 -923 256 -908
rect 254 -930 256 -927
rect 308 -952 310 -944
rect 308 -966 310 -960
rect 308 -984 310 -978
rect 308 -996 310 -992
rect 264 -1048 266 -1045
rect 308 -1052 310 -1045
rect 264 -1071 266 -1056
rect 308 -1066 310 -1060
rect 264 -1078 266 -1075
rect 308 -1084 310 -1078
rect 308 -1096 310 -1092
rect 308 -1162 310 -1155
rect 308 -1176 310 -1170
rect 308 -1194 310 -1188
rect 308 -1206 310 -1202
<< polycontact >>
rect 307 889 311 893
rect 307 835 311 839
rect 250 804 254 808
rect 307 780 311 784
rect 307 724 311 728
rect 307 679 311 683
rect 260 656 264 660
rect 307 624 311 628
rect 307 569 311 573
rect 307 514 311 518
rect 307 458 311 462
rect 307 404 311 408
rect 250 373 254 377
rect 307 349 311 353
rect 307 293 311 297
rect 307 248 311 252
rect 260 225 264 229
rect 307 193 311 197
rect 307 138 311 142
rect 307 83 311 87
rect 688 65 692 69
rect 731 65 735 69
rect 709 58 713 62
rect 851 39 855 43
rect 896 46 900 50
rect 913 42 917 46
rect 32 34 36 38
rect 12 17 16 21
rect 55 16 59 20
rect 75 13 79 17
rect 93 16 97 20
rect 130 16 134 20
rect 307 27 311 31
rect 870 20 874 24
rect 688 -10 692 -6
rect 731 -10 735 -6
rect 709 -17 713 -13
rect 32 -26 36 -22
rect 307 -27 311 -23
rect 12 -43 16 -39
rect 55 -44 59 -40
rect 75 -47 79 -43
rect 93 -44 97 -40
rect 130 -44 134 -40
rect 851 -39 855 -35
rect 896 -32 900 -28
rect 913 -36 917 -32
rect 250 -58 254 -54
rect 457 -68 461 -64
rect 500 -68 504 -64
rect 870 -58 874 -54
rect 479 -75 483 -71
rect 32 -86 36 -82
rect 307 -82 311 -78
rect 688 -85 692 -81
rect 731 -85 735 -81
rect 12 -103 16 -99
rect 55 -104 59 -100
rect 75 -107 79 -103
rect 93 -104 97 -100
rect 130 -104 134 -100
rect 709 -92 713 -88
rect 851 -117 855 -113
rect 896 -110 900 -106
rect 913 -114 917 -110
rect 468 -128 472 -124
rect 511 -128 515 -124
rect 307 -138 311 -134
rect 489 -135 493 -131
rect 870 -136 874 -132
rect 32 -146 36 -142
rect 12 -163 16 -159
rect 55 -164 59 -160
rect 75 -167 79 -163
rect 93 -164 97 -160
rect 130 -164 134 -160
rect 688 -160 692 -156
rect 731 -160 735 -156
rect 709 -167 713 -163
rect 307 -183 311 -179
rect 32 -206 36 -202
rect 260 -206 264 -202
rect 468 -188 472 -184
rect 511 -188 515 -184
rect 489 -195 493 -191
rect 851 -195 855 -191
rect 896 -188 900 -184
rect 913 -192 917 -188
rect 12 -223 16 -219
rect 55 -224 59 -220
rect 75 -227 79 -223
rect 93 -224 97 -220
rect 130 -224 134 -220
rect 870 -214 874 -210
rect 307 -238 311 -234
rect 468 -248 472 -244
rect 511 -248 515 -244
rect 489 -255 493 -251
rect 32 -276 36 -272
rect 851 -273 855 -269
rect 896 -266 900 -262
rect 913 -270 917 -266
rect 12 -293 16 -289
rect 55 -294 59 -290
rect 75 -297 79 -293
rect 93 -294 97 -290
rect 130 -294 134 -290
rect 307 -293 311 -289
rect 870 -292 874 -288
rect 468 -308 472 -304
rect 511 -308 515 -304
rect 489 -315 493 -311
rect 32 -336 36 -332
rect 12 -353 16 -349
rect 55 -354 59 -350
rect 75 -357 79 -353
rect 93 -354 97 -350
rect 130 -354 134 -350
rect 307 -348 311 -344
rect 32 -396 36 -392
rect 12 -413 16 -409
rect 55 -414 59 -410
rect 75 -417 79 -413
rect 93 -414 97 -410
rect 130 -414 134 -410
rect 307 -404 311 -400
rect 32 -456 36 -452
rect 307 -458 311 -454
rect 12 -473 16 -469
rect 55 -474 59 -470
rect 75 -477 79 -473
rect 93 -474 97 -470
rect 130 -474 134 -470
rect 250 -489 254 -485
rect 32 -516 36 -512
rect 307 -513 311 -509
rect 12 -533 16 -529
rect 55 -534 59 -530
rect 75 -537 79 -533
rect 93 -534 97 -530
rect 130 -534 134 -530
rect 307 -569 311 -565
rect 307 -614 311 -610
rect 260 -637 264 -633
rect 307 -669 311 -665
rect 307 -724 311 -720
rect 307 -779 311 -775
rect 307 -835 311 -831
rect 307 -889 311 -885
rect 250 -920 254 -916
rect 307 -944 311 -940
rect 307 -1000 311 -996
rect 307 -1045 311 -1041
rect 260 -1068 264 -1064
rect 307 -1100 311 -1096
rect 307 -1155 311 -1151
rect 307 -1210 311 -1206
<< metal1 >>
rect 307 893 311 896
rect 289 874 303 882
rect 315 874 329 882
rect 289 850 296 874
rect 315 859 319 866
rect 322 864 329 874
rect 322 850 329 857
rect 289 842 303 850
rect 315 842 329 850
rect 232 828 267 832
rect 232 684 236 828
rect 249 824 253 828
rect 257 808 261 816
rect 289 810 296 842
rect 272 808 296 810
rect 246 804 250 808
rect 257 804 296 808
rect 257 801 261 804
rect 272 803 296 804
rect 249 793 253 797
rect 246 789 267 793
rect 289 772 296 803
rect 307 800 311 835
rect 307 784 311 795
rect 289 764 303 772
rect 315 764 711 772
rect 289 740 296 764
rect 315 749 319 756
rect 322 740 329 764
rect 289 732 303 740
rect 315 732 329 740
rect 307 712 311 724
rect 268 710 271 711
rect 268 706 306 710
rect 232 680 277 684
rect 307 683 311 705
rect 232 401 236 680
rect 259 676 263 680
rect 322 678 329 732
rect 321 672 329 678
rect 267 660 271 668
rect 289 664 303 672
rect 315 664 329 672
rect 259 656 260 660
rect 267 656 276 660
rect 267 653 271 656
rect 259 645 263 649
rect 252 641 277 645
rect 289 640 296 664
rect 314 649 318 656
rect 321 653 329 664
rect 322 640 329 653
rect 289 632 303 640
rect 315 632 329 640
rect 289 599 296 632
rect 282 592 296 599
rect 289 562 296 592
rect 307 620 311 624
rect 307 573 311 615
rect 289 554 303 562
rect 315 554 329 562
rect 289 530 296 554
rect 315 539 319 546
rect 322 544 329 554
rect 322 530 329 537
rect 289 522 303 530
rect 315 522 329 530
rect 307 462 311 465
rect 289 443 303 451
rect 315 443 329 451
rect 289 419 296 443
rect 315 428 319 435
rect 322 433 329 443
rect 322 419 329 426
rect 289 411 303 419
rect 315 411 329 419
rect 232 397 267 401
rect 232 253 236 397
rect 249 393 253 397
rect 257 377 261 385
rect 289 379 296 411
rect 272 377 296 379
rect 246 373 250 377
rect 257 373 296 377
rect 257 370 261 373
rect 272 372 296 373
rect 249 362 253 366
rect 246 358 267 362
rect 289 341 296 372
rect 307 369 311 404
rect 307 353 311 364
rect 289 333 303 341
rect 315 333 611 341
rect 289 309 296 333
rect 315 318 319 325
rect 322 309 329 333
rect 289 301 303 309
rect 315 301 329 309
rect 307 281 311 293
rect 268 279 271 280
rect 268 275 306 279
rect 232 249 277 253
rect 307 252 311 274
rect 232 67 236 249
rect 259 245 263 249
rect 322 247 329 301
rect 321 241 329 247
rect 267 229 271 237
rect 289 233 303 241
rect 315 233 329 241
rect 259 225 260 229
rect 267 225 276 229
rect 267 222 271 225
rect 259 214 263 218
rect 252 210 277 214
rect 289 209 296 233
rect 314 218 318 225
rect 321 222 329 233
rect 322 209 329 222
rect 289 201 303 209
rect 315 201 329 209
rect 289 168 296 201
rect 282 161 296 168
rect 289 131 296 161
rect 307 189 311 193
rect 307 142 311 184
rect 596 146 604 333
rect 289 123 303 131
rect 315 123 329 131
rect 289 99 296 123
rect 315 108 319 115
rect 322 113 329 123
rect 638 124 646 764
rect 322 99 329 106
rect 289 91 303 99
rect 315 91 329 99
rect 527 94 679 95
rect 527 91 770 94
rect 232 63 455 67
rect 232 45 236 63
rect -8 41 236 45
rect -8 -15 -4 41
rect 9 34 13 41
rect 5 17 12 21
rect 25 13 29 26
rect 37 20 41 33
rect 52 34 56 41
rect 90 40 147 41
rect 90 34 94 40
rect 129 36 133 40
rect 64 26 82 30
rect 102 26 124 30
rect 37 16 55 20
rect 68 13 72 26
rect 78 23 82 26
rect 78 20 88 23
rect 21 9 37 13
rect 9 4 13 9
rect 84 16 93 20
rect 106 13 110 26
rect 121 20 124 26
rect 137 20 141 28
rect 121 16 130 20
rect 137 16 157 20
rect 137 13 141 16
rect 52 4 56 9
rect 90 5 94 9
rect 129 5 133 9
rect 90 4 142 5
rect 4 0 142 4
rect -8 -16 94 -15
rect -8 -19 147 -16
rect -8 -75 -4 -19
rect 9 -26 13 -19
rect 5 -43 12 -39
rect 25 -47 29 -34
rect 37 -40 41 -27
rect 52 -26 56 -19
rect 90 -20 147 -19
rect 90 -26 94 -20
rect 129 -24 133 -20
rect 64 -34 82 -30
rect 102 -34 124 -30
rect 37 -44 55 -40
rect 68 -47 72 -34
rect 78 -37 82 -34
rect 78 -40 88 -37
rect 21 -51 37 -47
rect 9 -56 13 -51
rect 84 -44 93 -40
rect 106 -47 110 -34
rect 121 -40 124 -34
rect 137 -40 141 -32
rect 190 -39 195 17
rect 150 -40 195 -39
rect 121 -44 130 -40
rect 137 -44 195 -40
rect 232 -30 236 41
rect 307 31 311 34
rect 289 12 303 20
rect 315 12 329 20
rect 289 -12 296 12
rect 315 -3 319 4
rect 322 2 329 12
rect 322 -12 329 -5
rect 289 -20 303 -12
rect 315 -20 329 -12
rect 232 -34 267 -30
rect 137 -47 141 -44
rect 52 -56 56 -51
rect 90 -55 94 -51
rect 129 -55 133 -51
rect 90 -56 147 -55
rect 4 -60 147 -56
rect -8 -76 94 -75
rect -8 -79 147 -76
rect -8 -135 -4 -79
rect 9 -86 13 -79
rect 5 -103 12 -99
rect 25 -107 29 -94
rect 37 -100 41 -87
rect 52 -86 56 -79
rect 90 -80 147 -79
rect 90 -86 94 -80
rect 129 -84 133 -80
rect 64 -94 82 -90
rect 102 -94 124 -90
rect 37 -104 55 -100
rect 68 -107 72 -94
rect 78 -97 82 -94
rect 78 -100 88 -97
rect 21 -111 37 -107
rect 9 -116 13 -111
rect 84 -104 93 -100
rect 106 -107 110 -94
rect 121 -100 124 -94
rect 137 -100 141 -92
rect 151 -97 185 -92
rect 151 -100 156 -97
rect 121 -104 130 -100
rect 137 -104 156 -100
rect 137 -107 141 -104
rect 52 -116 56 -111
rect 90 -115 94 -111
rect 129 -115 133 -111
rect 90 -116 147 -115
rect 4 -120 147 -116
rect -8 -136 94 -135
rect -8 -139 147 -136
rect -8 -195 -4 -139
rect 9 -146 13 -139
rect 5 -163 12 -159
rect 25 -167 29 -154
rect 37 -160 41 -147
rect 52 -146 56 -139
rect 90 -140 147 -139
rect 90 -146 94 -140
rect 129 -144 133 -140
rect 64 -154 82 -150
rect 102 -154 124 -150
rect 37 -164 55 -160
rect 68 -167 72 -154
rect 78 -157 82 -154
rect 78 -160 88 -157
rect 21 -171 37 -167
rect 9 -176 13 -171
rect 84 -164 93 -160
rect 106 -167 110 -154
rect 121 -160 124 -154
rect 137 -160 141 -152
rect 151 -160 156 -159
rect 121 -164 130 -160
rect 137 -162 156 -160
rect 137 -164 196 -162
rect 137 -167 141 -164
rect 151 -167 196 -164
rect 52 -176 56 -171
rect 90 -175 94 -171
rect 129 -175 133 -171
rect 90 -176 147 -175
rect 4 -180 147 -176
rect 232 -178 236 -34
rect 249 -38 253 -34
rect 257 -54 261 -46
rect 289 -52 296 -20
rect 272 -54 296 -52
rect 246 -58 250 -54
rect 257 -58 296 -54
rect 257 -61 261 -58
rect 272 -59 296 -58
rect 249 -69 253 -65
rect 246 -73 267 -69
rect 289 -90 296 -59
rect 307 -62 311 -27
rect 451 -39 455 63
rect 527 -39 531 91
rect 675 90 770 91
rect 689 85 693 90
rect 716 83 720 90
rect 732 83 736 90
rect 681 69 685 77
rect 724 69 728 75
rect 672 65 685 69
rect 692 65 728 69
rect 735 65 751 69
rect 681 62 685 65
rect 716 62 720 65
rect 678 58 681 62
rect 689 54 693 58
rect 626 53 700 54
rect 732 53 736 58
rect 626 49 738 53
rect 626 -17 631 49
rect 747 36 751 65
rect 708 31 747 35
rect 766 19 770 90
rect 675 15 770 19
rect 689 10 693 15
rect 716 8 720 15
rect 732 8 736 15
rect 681 -6 685 2
rect 724 -6 728 0
rect 672 -10 685 -6
rect 692 -10 728 -6
rect 735 -10 736 -6
rect 672 -11 676 -10
rect 668 -15 676 -11
rect 681 -13 685 -10
rect 716 -13 720 -10
rect 546 -21 631 -17
rect 689 -21 693 -17
rect 708 -17 709 -13
rect 625 -22 700 -21
rect 732 -22 736 -17
rect 625 -26 742 -22
rect 451 -43 532 -39
rect 456 -44 480 -43
rect 456 -50 460 -44
rect 472 -50 476 -44
rect 499 -46 503 -43
rect 464 -64 468 -58
rect 507 -64 511 -56
rect 307 -78 311 -67
rect 453 -68 457 -64
rect 464 -68 500 -64
rect 507 -68 514 -64
rect 472 -71 476 -68
rect 507 -71 511 -68
rect 483 -75 485 -71
rect 456 -80 460 -75
rect 499 -79 503 -75
rect 492 -80 509 -79
rect 450 -81 509 -80
rect 453 -84 509 -81
rect 289 -98 303 -90
rect 315 -98 427 -90
rect 289 -122 296 -98
rect 315 -113 319 -106
rect 322 -122 329 -98
rect 528 -99 532 -43
rect 572 -64 576 -34
rect 551 -68 577 -64
rect 626 -96 631 -26
rect 766 -56 770 15
rect 835 54 839 77
rect 850 73 954 77
rect 866 61 870 64
rect 835 49 836 54
rect 874 61 878 73
rect 882 61 886 64
rect 912 62 916 73
rect 835 31 839 49
rect 858 47 862 53
rect 896 50 900 54
rect 858 43 893 47
rect 920 46 924 54
rect 903 43 913 46
rect 849 39 851 43
rect 858 40 862 43
rect 882 40 886 43
rect 889 42 913 43
rect 920 42 937 46
rect 889 39 907 42
rect 920 39 924 42
rect 866 31 870 36
rect 912 31 916 35
rect 835 27 930 31
rect 675 -60 770 -56
rect 689 -65 693 -60
rect 716 -67 720 -60
rect 732 -67 736 -60
rect 681 -81 685 -73
rect 724 -81 728 -75
rect 674 -85 685 -81
rect 692 -85 728 -81
rect 735 -84 749 -81
rect 735 -85 743 -84
rect 674 -88 678 -85
rect 681 -88 685 -85
rect 716 -88 720 -85
rect 689 -96 693 -92
rect 708 -92 709 -88
rect 455 -103 532 -99
rect 625 -97 700 -96
rect 732 -97 736 -92
rect 625 -101 740 -97
rect 469 -108 473 -103
rect 289 -130 303 -122
rect 315 -130 329 -122
rect 496 -110 500 -103
rect 512 -110 516 -103
rect 461 -124 465 -116
rect 504 -124 508 -118
rect 528 -119 532 -103
rect 454 -127 465 -124
rect 307 -150 311 -138
rect 268 -152 271 -151
rect 268 -156 306 -152
rect 232 -182 277 -178
rect 307 -179 311 -157
rect -8 -196 94 -195
rect -8 -199 147 -196
rect -8 -265 -4 -199
rect 9 -206 13 -199
rect 5 -223 12 -219
rect 25 -227 29 -214
rect 37 -220 41 -207
rect 52 -206 56 -199
rect 90 -200 147 -199
rect 90 -206 94 -200
rect 129 -204 133 -200
rect 64 -214 82 -210
rect 102 -214 124 -210
rect 37 -224 55 -220
rect 68 -227 72 -214
rect 78 -217 82 -214
rect 78 -220 88 -217
rect 21 -231 37 -227
rect 9 -236 13 -231
rect 84 -224 93 -220
rect 106 -227 110 -214
rect 121 -220 124 -214
rect 137 -220 141 -212
rect 146 -220 185 -219
rect 121 -224 130 -220
rect 137 -224 185 -220
rect 137 -227 141 -224
rect 146 -225 185 -224
rect 52 -236 56 -231
rect 90 -235 94 -231
rect 129 -235 133 -231
rect 90 -236 147 -235
rect 4 -240 147 -236
rect -8 -266 94 -265
rect -8 -269 147 -266
rect -8 -325 -4 -269
rect 9 -276 13 -269
rect 5 -293 12 -289
rect 25 -297 29 -284
rect 37 -290 41 -277
rect 52 -276 56 -269
rect 90 -270 147 -269
rect 90 -276 94 -270
rect 129 -274 133 -270
rect 64 -284 82 -280
rect 102 -284 124 -280
rect 37 -294 55 -290
rect 68 -297 72 -284
rect 78 -287 82 -284
rect 78 -290 88 -287
rect 21 -301 37 -297
rect 9 -306 13 -301
rect 84 -294 93 -290
rect 106 -297 110 -284
rect 121 -290 124 -284
rect 137 -290 141 -282
rect 157 -290 160 -289
rect 121 -294 130 -290
rect 137 -294 160 -290
rect 137 -297 141 -294
rect 52 -306 56 -301
rect 90 -305 94 -301
rect 129 -305 133 -301
rect 90 -306 147 -305
rect 4 -310 147 -306
rect -8 -326 94 -325
rect -8 -329 147 -326
rect -8 -385 -4 -329
rect 9 -336 13 -329
rect 5 -353 12 -349
rect 25 -357 29 -344
rect 37 -350 41 -337
rect 52 -336 56 -329
rect 90 -330 147 -329
rect 90 -336 94 -330
rect 129 -334 133 -330
rect 64 -344 82 -340
rect 102 -344 124 -340
rect 37 -354 55 -350
rect 68 -357 72 -344
rect 78 -347 82 -344
rect 78 -350 88 -347
rect 21 -361 37 -357
rect 9 -366 13 -361
rect 84 -354 93 -350
rect 106 -357 110 -344
rect 121 -350 124 -344
rect 137 -350 141 -342
rect 206 -341 211 -306
rect 206 -350 211 -346
rect 121 -354 130 -350
rect 137 -354 211 -350
rect 137 -357 141 -354
rect 52 -366 56 -361
rect 90 -365 94 -361
rect 129 -365 133 -361
rect 90 -366 147 -365
rect 4 -370 147 -366
rect -8 -386 94 -385
rect -8 -389 147 -386
rect -8 -445 -4 -389
rect 9 -396 13 -389
rect 5 -413 12 -409
rect 25 -417 29 -404
rect 37 -410 41 -397
rect 52 -396 56 -389
rect 90 -390 147 -389
rect 90 -396 94 -390
rect 129 -394 133 -390
rect 64 -404 82 -400
rect 102 -404 124 -400
rect 37 -414 55 -410
rect 68 -417 72 -404
rect 78 -407 82 -404
rect 78 -410 88 -407
rect 21 -421 37 -417
rect 9 -426 13 -421
rect 84 -414 93 -410
rect 106 -417 110 -404
rect 121 -410 124 -404
rect 137 -410 141 -402
rect 154 -410 159 -409
rect 121 -414 130 -410
rect 137 -414 159 -410
rect 137 -417 141 -414
rect 52 -426 56 -421
rect 154 -419 159 -414
rect 90 -425 94 -421
rect 129 -425 133 -421
rect 90 -426 147 -425
rect 4 -430 147 -426
rect -8 -446 94 -445
rect -8 -449 147 -446
rect -8 -505 -4 -449
rect 9 -456 13 -449
rect 5 -473 12 -469
rect 25 -477 29 -464
rect 37 -470 41 -457
rect 52 -456 56 -449
rect 90 -450 147 -449
rect 90 -456 94 -450
rect 129 -454 133 -450
rect 64 -464 82 -460
rect 102 -464 124 -460
rect 37 -474 55 -470
rect 68 -477 72 -464
rect 78 -467 82 -464
rect 78 -470 88 -467
rect 21 -481 37 -477
rect 9 -486 13 -481
rect 84 -474 93 -470
rect 106 -477 110 -464
rect 121 -470 124 -464
rect 137 -470 141 -462
rect 232 -461 236 -182
rect 259 -186 263 -182
rect 322 -184 329 -130
rect 458 -128 465 -127
rect 472 -128 508 -124
rect 515 -128 521 -124
rect 461 -131 465 -128
rect 496 -131 500 -128
rect 529 -130 533 -119
rect 469 -139 473 -135
rect 488 -135 489 -131
rect 455 -140 480 -139
rect 512 -140 516 -135
rect 460 -144 522 -140
rect 321 -190 329 -184
rect 446 -155 516 -151
rect 446 -184 450 -155
rect 528 -159 532 -130
rect 455 -163 532 -159
rect 469 -168 473 -163
rect 496 -170 500 -163
rect 512 -170 516 -163
rect 461 -184 465 -176
rect 504 -184 508 -178
rect 267 -202 271 -194
rect 289 -198 303 -190
rect 315 -198 329 -190
rect 259 -206 260 -202
rect 267 -206 276 -202
rect 267 -209 271 -206
rect 259 -217 263 -213
rect 252 -221 277 -217
rect 289 -222 296 -198
rect 314 -213 318 -206
rect 321 -209 329 -198
rect 322 -222 329 -209
rect 289 -230 303 -222
rect 315 -230 329 -222
rect 446 -188 465 -184
rect 472 -187 508 -184
rect 472 -188 481 -187
rect 492 -188 508 -187
rect 515 -188 518 -184
rect 289 -263 296 -230
rect 282 -270 296 -263
rect 289 -300 296 -270
rect 307 -242 311 -238
rect 307 -289 311 -247
rect 372 -263 378 -192
rect 461 -191 465 -188
rect 496 -191 500 -188
rect 451 -199 457 -198
rect 469 -199 473 -195
rect 451 -200 480 -199
rect 512 -200 516 -195
rect 451 -203 522 -200
rect 455 -204 522 -203
rect 446 -214 519 -210
rect 446 -244 450 -214
rect 528 -219 532 -163
rect 455 -223 532 -219
rect 469 -228 473 -223
rect 496 -230 500 -223
rect 512 -230 516 -223
rect 461 -244 465 -236
rect 504 -244 508 -238
rect 401 -249 437 -244
rect 446 -248 465 -244
rect 472 -248 508 -244
rect 515 -248 517 -244
rect 323 -269 379 -263
rect 289 -308 303 -300
rect 315 -308 329 -300
rect 289 -332 296 -308
rect 315 -323 319 -316
rect 322 -318 329 -308
rect 322 -332 329 -325
rect 289 -340 303 -332
rect 315 -340 329 -332
rect 307 -400 311 -397
rect 289 -419 303 -411
rect 315 -419 329 -411
rect 289 -443 296 -419
rect 315 -434 319 -427
rect 322 -429 329 -419
rect 322 -443 329 -436
rect 289 -451 303 -443
rect 315 -451 329 -443
rect 232 -465 267 -461
rect 153 -470 159 -469
rect 121 -474 130 -470
rect 137 -474 159 -470
rect 137 -477 141 -474
rect 52 -486 56 -481
rect 90 -485 94 -481
rect 129 -485 133 -481
rect 90 -486 147 -485
rect 4 -490 147 -486
rect -8 -506 94 -505
rect -8 -509 147 -506
rect 9 -516 13 -509
rect 5 -533 12 -529
rect 25 -537 29 -524
rect 37 -530 41 -517
rect 52 -516 56 -509
rect 90 -510 147 -509
rect 90 -516 94 -510
rect 129 -514 133 -510
rect 64 -524 82 -520
rect 102 -524 124 -520
rect 37 -534 55 -530
rect 68 -537 72 -524
rect 78 -527 82 -524
rect 78 -530 88 -527
rect 21 -541 37 -537
rect 9 -546 13 -541
rect 84 -534 93 -530
rect 106 -537 110 -524
rect 121 -530 124 -524
rect 137 -530 141 -522
rect 152 -530 157 -529
rect 121 -534 130 -530
rect 137 -532 157 -530
rect 137 -534 172 -532
rect 137 -537 141 -534
rect 152 -537 172 -534
rect 52 -546 56 -541
rect 90 -545 94 -541
rect 129 -545 133 -541
rect 90 -546 147 -545
rect 4 -550 147 -546
rect 232 -609 236 -465
rect 249 -469 253 -465
rect 257 -485 261 -477
rect 289 -483 296 -451
rect 272 -485 296 -483
rect 246 -489 250 -485
rect 257 -489 296 -485
rect 257 -492 261 -489
rect 272 -490 296 -489
rect 249 -500 253 -496
rect 246 -504 267 -500
rect 289 -521 296 -490
rect 307 -493 311 -458
rect 307 -509 311 -498
rect 401 -502 406 -249
rect 432 -269 437 -249
rect 461 -251 465 -248
rect 496 -251 500 -248
rect 469 -259 473 -255
rect 488 -255 489 -251
rect 452 -260 480 -259
rect 512 -260 516 -255
rect 452 -263 522 -260
rect 447 -264 522 -263
rect 432 -274 517 -269
rect 528 -279 532 -223
rect 455 -283 532 -279
rect 469 -288 473 -283
rect 496 -290 500 -283
rect 512 -290 516 -283
rect 461 -304 465 -296
rect 504 -304 508 -298
rect 415 -308 465 -304
rect 472 -308 508 -304
rect 515 -308 533 -304
rect 415 -414 419 -308
rect 461 -311 465 -308
rect 496 -311 500 -308
rect 461 -316 465 -315
rect 469 -319 473 -315
rect 487 -315 489 -311
rect 451 -320 480 -319
rect 512 -320 516 -315
rect 451 -324 522 -320
rect 527 -338 533 -308
rect 433 -344 533 -338
rect 433 -353 439 -344
rect 415 -418 580 -414
rect 328 -507 406 -502
rect 598 -521 606 -125
rect 626 -171 631 -101
rect 745 -124 749 -106
rect 709 -128 749 -124
rect 766 -131 770 -60
rect 820 -67 824 -39
rect 835 -47 839 27
rect 867 20 870 24
rect 933 11 937 42
rect 950 -1 954 73
rect 852 -5 954 -1
rect 866 -17 870 -14
rect 874 -17 878 -5
rect 882 -17 886 -14
rect 912 -16 916 -5
rect 858 -31 862 -25
rect 896 -28 900 -24
rect 858 -35 893 -31
rect 920 -32 924 -24
rect 903 -35 913 -32
rect 848 -39 851 -35
rect 858 -38 862 -35
rect 882 -38 886 -35
rect 889 -36 913 -35
rect 920 -36 937 -32
rect 889 -39 907 -36
rect 920 -39 924 -36
rect 866 -47 870 -42
rect 912 -47 916 -43
rect 835 -51 930 -47
rect 675 -135 770 -131
rect 835 -125 839 -51
rect 866 -58 870 -54
rect 845 -113 849 -60
rect 933 -68 937 -36
rect 950 -79 954 -5
rect 852 -83 954 -79
rect 866 -95 870 -92
rect 874 -95 878 -83
rect 882 -95 886 -92
rect 912 -94 916 -83
rect 858 -109 862 -103
rect 896 -106 900 -102
rect 858 -113 893 -109
rect 920 -110 924 -102
rect 903 -113 913 -110
rect 845 -117 851 -113
rect 858 -116 862 -113
rect 882 -116 886 -113
rect 889 -114 913 -113
rect 920 -114 933 -110
rect 889 -117 907 -114
rect 920 -117 924 -114
rect 866 -125 870 -120
rect 912 -125 916 -121
rect 835 -129 930 -125
rect 689 -140 693 -135
rect 716 -142 720 -135
rect 732 -142 736 -135
rect 681 -156 685 -148
rect 724 -156 728 -150
rect 678 -160 685 -156
rect 692 -160 728 -156
rect 681 -163 685 -160
rect 716 -163 720 -160
rect 689 -171 693 -167
rect 626 -172 700 -171
rect 732 -172 736 -167
rect 626 -176 742 -172
rect 835 -203 839 -129
rect 867 -136 870 -132
rect 950 -157 954 -83
rect 852 -161 954 -157
rect 866 -173 870 -170
rect 874 -173 878 -161
rect 882 -173 886 -170
rect 912 -172 916 -161
rect 858 -187 862 -181
rect 858 -191 893 -187
rect 920 -188 924 -180
rect 903 -191 913 -188
rect 849 -195 851 -191
rect 858 -194 862 -191
rect 882 -194 886 -191
rect 889 -192 913 -191
rect 920 -192 937 -188
rect 889 -195 907 -192
rect 920 -195 924 -192
rect 866 -203 870 -198
rect 912 -203 916 -199
rect 835 -207 930 -203
rect 835 -281 839 -207
rect 865 -214 870 -210
rect 933 -225 937 -192
rect 950 -235 954 -161
rect 852 -239 954 -235
rect 866 -251 870 -248
rect 874 -251 878 -239
rect 882 -251 886 -248
rect 912 -250 916 -239
rect 858 -265 862 -259
rect 896 -260 898 -256
rect 896 -262 900 -260
rect 858 -269 893 -265
rect 920 -266 924 -258
rect 903 -269 913 -266
rect 849 -273 851 -269
rect 858 -272 862 -269
rect 882 -272 886 -269
rect 889 -270 913 -269
rect 920 -270 933 -266
rect 889 -273 907 -270
rect 920 -273 924 -270
rect 866 -281 870 -276
rect 912 -281 916 -277
rect 835 -285 930 -281
rect 863 -292 870 -288
rect 874 -292 933 -288
rect 904 -331 943 -327
rect 896 -335 943 -331
rect 289 -529 303 -521
rect 315 -529 606 -521
rect 289 -553 296 -529
rect 315 -544 319 -537
rect 322 -553 329 -529
rect 289 -561 303 -553
rect 315 -561 329 -553
rect 307 -581 311 -569
rect 268 -583 271 -582
rect 268 -587 306 -583
rect 232 -613 277 -609
rect 307 -610 311 -588
rect 232 -892 236 -613
rect 259 -617 263 -613
rect 322 -615 329 -561
rect 321 -621 329 -615
rect 267 -633 271 -625
rect 289 -629 303 -621
rect 315 -629 329 -621
rect 259 -637 260 -633
rect 267 -637 276 -633
rect 267 -640 271 -637
rect 259 -648 263 -644
rect 252 -652 277 -648
rect 289 -653 296 -629
rect 314 -644 318 -637
rect 321 -640 329 -629
rect 322 -653 329 -640
rect 289 -661 303 -653
rect 315 -661 329 -653
rect 289 -694 296 -661
rect 282 -701 296 -694
rect 289 -731 296 -701
rect 307 -673 311 -669
rect 307 -720 311 -678
rect 289 -739 303 -731
rect 315 -739 329 -731
rect 289 -763 296 -739
rect 315 -754 319 -747
rect 322 -749 329 -739
rect 322 -763 329 -756
rect 289 -771 303 -763
rect 315 -771 329 -763
rect 307 -831 311 -828
rect 289 -850 303 -842
rect 315 -850 329 -842
rect 289 -874 296 -850
rect 315 -865 319 -858
rect 322 -860 329 -850
rect 322 -874 329 -867
rect 289 -882 303 -874
rect 315 -882 329 -874
rect 232 -896 267 -892
rect 232 -1040 236 -896
rect 249 -900 253 -896
rect 257 -916 261 -908
rect 289 -914 296 -882
rect 272 -916 296 -914
rect 246 -920 250 -916
rect 257 -920 296 -916
rect 257 -923 261 -920
rect 272 -921 296 -920
rect 249 -931 253 -927
rect 246 -935 267 -931
rect 289 -952 296 -921
rect 307 -924 311 -889
rect 307 -940 311 -929
rect 935 -952 943 -335
rect 289 -960 303 -952
rect 315 -960 943 -952
rect 289 -984 296 -960
rect 315 -975 319 -968
rect 322 -984 329 -960
rect 289 -992 303 -984
rect 315 -992 329 -984
rect 307 -1012 311 -1000
rect 268 -1014 271 -1013
rect 268 -1018 306 -1014
rect 232 -1044 277 -1040
rect 307 -1041 311 -1019
rect 259 -1048 263 -1044
rect 322 -1046 329 -992
rect 321 -1052 329 -1046
rect 267 -1064 271 -1056
rect 289 -1060 303 -1052
rect 315 -1060 329 -1052
rect 259 -1068 260 -1064
rect 267 -1068 276 -1064
rect 267 -1071 271 -1068
rect 259 -1079 263 -1075
rect 252 -1083 277 -1079
rect 289 -1084 296 -1060
rect 314 -1075 318 -1068
rect 321 -1071 329 -1060
rect 322 -1084 329 -1071
rect 289 -1092 303 -1084
rect 315 -1092 329 -1084
rect 289 -1125 296 -1092
rect 282 -1132 296 -1125
rect 289 -1162 296 -1132
rect 307 -1104 311 -1100
rect 307 -1151 311 -1109
rect 289 -1170 303 -1162
rect 315 -1170 329 -1162
rect 289 -1194 296 -1170
rect 315 -1185 319 -1178
rect 322 -1180 329 -1170
rect 322 -1194 329 -1187
rect 289 -1202 303 -1194
rect 315 -1202 329 -1194
<< m2contact >>
rect 322 857 329 864
rect 241 788 246 793
rect 307 795 312 800
rect 276 656 281 661
rect 247 640 252 645
rect 307 615 312 620
rect 322 537 329 544
rect 322 426 329 433
rect 241 357 246 362
rect 307 364 312 369
rect 611 333 619 341
rect 276 225 281 230
rect 247 209 252 214
rect 307 184 312 189
rect 596 138 604 146
rect 638 116 646 124
rect 322 106 329 113
rect 36 33 41 38
rect -1 0 4 5
rect 37 8 42 13
rect 152 20 157 25
rect 190 17 195 22
rect 75 8 80 13
rect 142 0 147 5
rect 36 -27 41 -22
rect -1 -60 4 -55
rect 37 -52 42 -47
rect 322 -5 329 2
rect 75 -52 80 -47
rect 36 -87 41 -82
rect -1 -120 4 -115
rect 37 -112 42 -107
rect 185 -97 190 -92
rect 75 -112 80 -107
rect 36 -147 41 -142
rect -1 -180 4 -175
rect 37 -172 42 -167
rect 196 -167 201 -162
rect 75 -172 80 -167
rect 241 -74 246 -69
rect 673 57 678 62
rect 704 57 709 62
rect 540 -22 546 -16
rect 738 48 743 53
rect 703 31 708 36
rect 747 31 752 36
rect 703 -18 708 -13
rect 572 -34 577 -29
rect 307 -67 312 -62
rect 514 -68 519 -63
rect 448 -86 453 -81
rect 546 -68 551 -63
rect 866 64 871 69
rect 836 49 841 54
rect 882 64 887 69
rect 896 54 901 59
rect 844 39 849 44
rect 673 -93 678 -88
rect 703 -93 708 -88
rect 36 -207 41 -202
rect -1 -240 4 -235
rect 37 -232 42 -227
rect 185 -225 191 -219
rect 75 -232 80 -227
rect 36 -277 41 -272
rect -1 -310 4 -305
rect 37 -302 42 -297
rect 75 -302 80 -297
rect 36 -337 41 -332
rect -1 -370 4 -365
rect 37 -362 42 -357
rect 75 -362 80 -357
rect 36 -397 41 -392
rect -1 -430 4 -425
rect 37 -422 42 -417
rect 75 -422 80 -417
rect 36 -457 41 -452
rect -1 -490 4 -485
rect 37 -482 42 -477
rect 598 -125 606 -117
rect 483 -136 488 -131
rect 455 -145 460 -140
rect 516 -155 521 -150
rect 276 -206 281 -201
rect 247 -222 252 -217
rect 307 -247 312 -242
rect 446 -203 451 -198
rect 519 -214 524 -209
rect 517 -248 522 -243
rect 322 -325 329 -318
rect 322 -436 329 -429
rect 75 -482 80 -477
rect 36 -517 41 -512
rect -1 -550 4 -545
rect 37 -542 42 -537
rect 75 -542 80 -537
rect 241 -505 246 -500
rect 307 -498 312 -493
rect 447 -263 452 -258
rect 517 -274 522 -269
rect 446 -324 451 -319
rect 433 -359 439 -353
rect 580 -418 585 -413
rect 323 -507 328 -502
rect 704 -128 709 -123
rect 820 -39 825 -34
rect 862 19 867 24
rect 933 6 938 11
rect 866 -14 871 -9
rect 882 -14 887 -9
rect 843 -39 848 -34
rect 820 -72 825 -67
rect 845 -60 850 -55
rect 860 -60 866 -54
rect 933 -73 938 -68
rect 866 -92 871 -87
rect 882 -92 887 -87
rect 673 -160 678 -155
rect 735 -160 740 -155
rect 704 -168 709 -163
rect 862 -137 867 -132
rect 866 -170 871 -165
rect 882 -170 887 -165
rect 896 -184 901 -179
rect 844 -196 849 -191
rect 933 -230 938 -225
rect 866 -248 871 -243
rect 882 -248 887 -243
rect 898 -260 903 -255
rect 844 -274 849 -269
rect 933 -292 938 -287
rect 896 -331 904 -324
rect 276 -637 281 -632
rect 247 -653 252 -648
rect 307 -678 312 -673
rect 322 -756 329 -749
rect 322 -867 329 -860
rect 241 -936 246 -931
rect 307 -929 312 -924
rect 276 -1068 281 -1063
rect 247 -1084 252 -1079
rect 307 -1109 312 -1104
rect 322 -1187 329 -1180
<< pm12contact >>
rect 113 15 118 20
rect 113 -45 118 -40
rect 113 -105 118 -100
rect 113 -165 118 -160
rect 113 -225 118 -220
rect 113 -295 118 -290
rect 113 -355 118 -350
rect 113 -415 118 -410
rect 113 -475 118 -470
rect 113 -535 118 -530
<< metal2 >>
rect 329 857 346 864
rect 281 795 307 799
rect 151 706 224 711
rect 151 705 203 706
rect 151 96 157 705
rect 242 645 246 788
rect 242 640 247 645
rect 242 388 246 640
rect 281 619 285 795
rect 339 650 346 857
rect 339 643 362 650
rect 281 615 307 619
rect 339 544 346 643
rect 329 537 346 544
rect 380 479 381 484
rect 329 426 346 433
rect 237 384 246 388
rect 237 382 242 384
rect 237 376 241 382
rect 234 373 241 376
rect 237 369 241 373
rect 237 365 246 369
rect 241 362 246 365
rect 37 48 117 52
rect 37 38 41 48
rect 113 20 117 48
rect 152 25 157 96
rect 190 281 195 282
rect 190 280 221 281
rect 190 276 224 280
rect 190 22 195 276
rect 212 275 224 276
rect 242 214 246 357
rect 281 364 307 368
rect 242 209 247 214
rect 242 58 246 209
rect 281 188 285 364
rect 339 219 346 426
rect 380 286 386 479
rect 619 333 897 341
rect 352 280 386 286
rect 352 245 358 280
rect 373 253 561 257
rect 352 239 388 245
rect 339 212 362 219
rect 281 184 307 188
rect 339 113 346 212
rect 329 106 346 113
rect 382 86 388 239
rect 242 54 444 58
rect 42 8 75 13
rect 242 5 246 54
rect 147 0 247 5
rect -1 -55 3 0
rect 37 -12 117 -8
rect 37 -22 41 -12
rect 113 -40 117 -12
rect 242 -43 246 0
rect 329 -5 346 2
rect 237 -47 246 -43
rect 42 -52 75 -47
rect 237 -49 242 -47
rect 237 -55 241 -49
rect 234 -58 241 -55
rect -1 -115 3 -60
rect 237 -62 241 -58
rect 237 -66 246 -62
rect 37 -72 117 -68
rect 37 -82 41 -72
rect 113 -100 117 -72
rect 241 -69 246 -66
rect 42 -112 75 -107
rect -1 -175 3 -120
rect 37 -132 117 -128
rect 37 -142 41 -132
rect 113 -160 117 -132
rect 185 -151 190 -97
rect 185 -156 224 -151
rect 42 -172 75 -167
rect -1 -235 3 -180
rect 37 -192 117 -188
rect 37 -202 41 -192
rect 113 -220 117 -192
rect 42 -232 75 -227
rect -1 -305 3 -240
rect 37 -262 117 -258
rect 37 -272 41 -262
rect 113 -290 117 -262
rect 42 -302 75 -297
rect -1 -365 3 -310
rect 37 -322 117 -318
rect 37 -332 41 -322
rect 113 -350 117 -322
rect 42 -362 75 -357
rect -1 -425 3 -370
rect 37 -382 117 -378
rect 37 -392 41 -382
rect 113 -410 117 -382
rect 42 -422 75 -417
rect -1 -485 3 -430
rect 37 -442 117 -438
rect 37 -452 41 -442
rect 113 -470 117 -442
rect 42 -482 75 -477
rect -1 -545 3 -490
rect 37 -502 117 -498
rect 37 -512 41 -502
rect 113 -530 117 -502
rect 42 -542 75 -537
rect 185 -1013 191 -225
rect 196 -582 201 -167
rect 242 -217 246 -74
rect 281 -67 307 -63
rect 242 -223 247 -217
rect 242 -474 246 -223
rect 281 -243 285 -67
rect 339 -212 346 -5
rect 440 -17 444 54
rect 440 -21 540 -17
rect 440 -81 444 -21
rect 519 -68 546 -64
rect 440 -85 448 -81
rect 440 -141 444 -85
rect 557 -131 561 253
rect 604 145 705 146
rect 604 138 709 145
rect 638 62 646 116
rect 703 62 709 138
rect 889 106 897 333
rect 889 100 900 106
rect 871 64 882 68
rect 638 57 673 62
rect 703 57 704 62
rect 896 59 900 100
rect 743 49 836 53
rect 572 40 830 44
rect 572 -29 576 40
rect 703 -13 707 31
rect 568 -107 573 -49
rect 747 -75 751 31
rect 826 24 830 40
rect 826 20 862 24
rect 810 -20 815 14
rect 871 -14 882 -10
rect 810 -25 846 -20
rect 851 -25 852 -20
rect 933 -20 937 6
rect 933 -24 946 -20
rect 792 -39 795 -32
rect 825 -39 843 -35
rect 756 -40 813 -39
rect 756 -45 757 -40
rect 762 -44 813 -40
rect 762 -45 825 -44
rect 747 -79 758 -75
rect 674 -102 678 -93
rect 674 -106 688 -102
rect 703 -110 708 -93
rect 643 -117 725 -110
rect 606 -118 725 -117
rect 606 -125 651 -118
rect 488 -135 561 -131
rect 440 -145 455 -141
rect 460 -145 462 -141
rect 440 -198 444 -145
rect 521 -155 578 -151
rect 573 -186 577 -155
rect 673 -172 677 -160
rect 704 -163 708 -128
rect 754 -156 758 -79
rect 740 -160 758 -156
rect 673 -176 758 -172
rect 792 -173 795 -45
rect 807 -50 825 -45
rect 803 -59 845 -55
rect 803 -186 807 -59
rect 850 -59 860 -55
rect 573 -190 807 -186
rect 440 -203 446 -198
rect 339 -219 362 -212
rect 281 -247 307 -243
rect 339 -318 346 -219
rect 329 -325 346 -318
rect 440 -258 444 -203
rect 820 -210 824 -72
rect 843 -76 906 -71
rect 843 -131 848 -76
rect 871 -92 882 -88
rect 843 -136 862 -131
rect 933 -144 937 -73
rect 845 -148 937 -144
rect 845 -191 849 -148
rect 942 -162 946 -24
rect 871 -170 882 -166
rect 896 -166 946 -162
rect 896 -179 900 -166
rect 524 -214 824 -210
rect 871 -248 882 -244
rect 440 -263 447 -258
rect 440 -266 445 -263
rect 440 -319 444 -266
rect 517 -269 522 -248
rect 619 -278 849 -274
rect 440 -324 446 -319
rect 439 -359 466 -353
rect 329 -436 346 -429
rect 237 -478 246 -474
rect 237 -480 242 -478
rect 237 -486 241 -480
rect 234 -489 241 -486
rect 237 -493 241 -489
rect 237 -497 246 -493
rect 241 -500 246 -497
rect 196 -587 224 -582
rect 242 -648 246 -505
rect 281 -498 307 -494
rect 242 -653 247 -648
rect 242 -905 246 -653
rect 281 -674 285 -498
rect 293 -567 299 -566
rect 293 -572 294 -567
rect 323 -572 328 -507
rect 293 -577 328 -572
rect 339 -643 346 -436
rect 339 -650 362 -643
rect 281 -678 307 -674
rect 339 -749 346 -650
rect 329 -756 346 -749
rect 460 -755 466 -359
rect 619 -414 623 -278
rect 898 -324 902 -260
rect 933 -287 937 -230
rect 933 -293 937 -292
rect 585 -418 623 -414
rect 378 -756 466 -755
rect 378 -761 379 -756
rect 384 -761 466 -756
rect 329 -867 346 -860
rect 237 -909 246 -905
rect 237 -911 242 -909
rect 237 -917 241 -911
rect 234 -920 241 -917
rect 237 -924 241 -920
rect 237 -928 246 -924
rect 241 -931 246 -928
rect 185 -1018 224 -1013
rect 185 -1019 202 -1018
rect 242 -1079 246 -936
rect 281 -929 307 -925
rect 242 -1083 247 -1079
rect 281 -1105 285 -929
rect 339 -1074 346 -867
rect 339 -1081 362 -1074
rect 281 -1109 307 -1105
rect 339 -1180 346 -1081
rect 329 -1187 346 -1180
<< m3contact >>
rect 224 706 229 711
rect 381 479 386 484
rect 245 373 250 378
rect 224 275 229 280
rect 368 253 373 258
rect 382 81 388 86
rect 245 -58 250 -53
rect 224 -156 229 -151
rect 568 -49 573 -44
rect 810 14 815 19
rect 846 -25 851 -20
rect 789 -32 796 -25
rect 757 -45 762 -40
rect 688 -106 693 -101
rect 568 -112 573 -107
rect 725 -118 731 -110
rect 825 -50 830 -44
rect 791 -178 796 -173
rect 906 -76 911 -71
rect 245 -489 250 -484
rect 224 -587 229 -582
rect 294 -572 299 -567
rect 379 -761 384 -756
rect 245 -920 250 -915
rect 224 -1018 229 -1013
<< m123contact >>
rect 306 896 313 903
rect 239 803 246 810
rect 263 706 268 711
rect 252 656 259 663
rect 306 705 313 712
rect 271 591 282 600
rect 306 507 313 514
rect 306 465 313 472
rect 263 275 268 280
rect 252 225 259 232
rect 306 274 313 281
rect 271 160 282 169
rect 306 76 313 83
rect 306 34 313 41
rect 160 -294 165 -289
rect 159 -419 164 -414
rect 159 -474 164 -469
rect 172 -537 177 -532
rect 263 -156 268 -151
rect 252 -206 259 -199
rect 206 -346 211 -341
rect 306 -157 313 -150
rect 448 -69 453 -64
rect 485 -76 490 -71
rect 427 -98 435 -90
rect 521 -127 526 -122
rect 453 -132 458 -127
rect 736 -10 742 -4
rect 844 39 849 44
rect 896 -24 901 -19
rect 743 -90 749 -84
rect 743 -106 750 -99
rect 372 -192 378 -186
rect 518 -188 523 -183
rect 484 -195 489 -190
rect 271 -271 282 -262
rect 316 -270 323 -263
rect 896 -102 901 -96
rect 860 -215 865 -210
rect 483 -256 488 -251
rect 482 -316 487 -311
rect 306 -355 313 -348
rect 306 -397 313 -390
rect 263 -587 268 -582
rect 252 -637 259 -630
rect 306 -588 313 -581
rect 271 -702 282 -693
rect 306 -786 313 -779
rect 306 -828 313 -821
rect 263 -1018 268 -1013
rect 252 -1068 259 -1061
rect 306 -1019 313 -1012
rect 271 -1133 282 -1124
rect 306 -1217 313 -1210
<< metal3 >>
rect 313 897 336 901
rect 212 804 239 808
rect 212 598 218 804
rect 223 711 230 712
rect 262 711 269 712
rect 223 706 224 711
rect 229 706 263 711
rect 268 706 269 711
rect 223 705 230 706
rect 252 663 256 706
rect 262 705 269 706
rect 332 710 336 897
rect 313 706 336 710
rect 332 676 336 706
rect 332 672 499 676
rect 251 656 252 662
rect 251 655 258 656
rect 167 593 271 598
rect 167 -284 172 593
rect 212 592 271 593
rect 260 501 266 592
rect 332 512 336 672
rect 313 508 336 512
rect 260 495 409 501
rect 380 484 387 485
rect 212 479 381 484
rect 386 479 387 484
rect 212 478 387 479
rect 212 377 218 478
rect 313 466 336 470
rect 244 378 251 379
rect 234 377 245 378
rect 212 373 245 377
rect 250 373 251 378
rect 212 172 218 373
rect 244 372 251 373
rect 223 280 230 281
rect 262 280 269 281
rect 223 275 224 280
rect 229 275 263 280
rect 268 275 269 280
rect 223 274 230 275
rect 252 232 256 275
rect 262 274 269 275
rect 332 279 336 466
rect 313 275 336 279
rect 332 257 336 275
rect 367 258 374 259
rect 367 257 368 258
rect 332 253 368 257
rect 373 253 374 258
rect 251 225 252 231
rect 251 224 258 225
rect 166 -288 172 -284
rect 159 -289 172 -288
rect 159 -294 160 -289
rect 165 -294 172 -289
rect 201 167 218 172
rect 159 -295 166 -294
rect 201 -295 206 167
rect 212 161 271 167
rect 332 81 336 253
rect 367 252 374 253
rect 313 77 336 81
rect 381 86 389 87
rect 381 81 382 86
rect 388 81 389 86
rect 381 80 389 81
rect 313 35 336 39
rect 244 -53 251 -52
rect 234 -54 245 -53
rect 212 -58 245 -54
rect 250 -58 251 -53
rect 212 -262 218 -58
rect 244 -59 251 -58
rect 223 -151 230 -150
rect 262 -151 269 -150
rect 223 -156 224 -151
rect 229 -156 263 -151
rect 268 -156 269 -151
rect 223 -157 230 -156
rect 252 -199 256 -156
rect 262 -157 269 -156
rect 332 -152 336 35
rect 382 -124 388 80
rect 403 -63 409 495
rect 495 -23 499 672
rect 485 -27 499 -23
rect 568 46 573 47
rect 568 44 849 46
rect 568 41 844 44
rect 403 -69 448 -63
rect 485 -70 489 -27
rect 568 -43 573 41
rect 809 19 816 20
rect 809 14 810 19
rect 815 18 816 19
rect 830 18 835 41
rect 815 14 835 18
rect 809 13 835 14
rect 800 3 900 9
rect 736 -4 742 -3
rect 595 -6 603 -5
rect 595 -12 661 -6
rect 567 -44 574 -43
rect 567 -49 568 -44
rect 573 -49 574 -44
rect 567 -50 574 -49
rect 484 -71 491 -70
rect 484 -76 485 -71
rect 490 -76 491 -71
rect 484 -77 491 -76
rect 426 -90 436 -89
rect 595 -90 603 -12
rect 655 -28 661 -12
rect 736 -28 742 -10
rect 655 -34 745 -28
rect 773 -30 789 -27
rect 655 -40 661 -34
rect 756 -40 763 -39
rect 655 -45 757 -40
rect 762 -45 763 -40
rect 655 -46 763 -45
rect 746 -81 752 -46
rect 745 -84 752 -81
rect 749 -89 752 -84
rect 426 -98 427 -90
rect 435 -98 603 -90
rect 426 -99 436 -98
rect 687 -101 694 -100
rect 687 -106 688 -101
rect 693 -105 743 -101
rect 693 -106 694 -105
rect 773 -101 776 -30
rect 750 -105 776 -101
rect 780 -39 788 -38
rect 800 -39 806 3
rect 896 -19 900 3
rect 845 -20 852 -19
rect 845 -25 846 -20
rect 851 -25 852 -20
rect 845 -26 852 -25
rect 780 -45 806 -39
rect 824 -44 831 -43
rect 567 -107 574 -106
rect 687 -107 694 -106
rect 567 -112 568 -107
rect 573 -112 574 -107
rect 567 -113 574 -112
rect 724 -110 732 -109
rect 780 -110 788 -45
rect 824 -50 825 -44
rect 830 -50 831 -44
rect 824 -51 831 -50
rect 846 -48 851 -26
rect 824 -63 830 -51
rect 846 -53 911 -48
rect 824 -69 901 -63
rect 896 -96 901 -69
rect 906 -70 911 -53
rect 905 -71 912 -70
rect 905 -76 906 -71
rect 911 -76 912 -71
rect 905 -77 912 -76
rect 445 -122 524 -117
rect 445 -124 449 -122
rect 382 -130 449 -124
rect 458 -132 463 -130
rect 453 -135 463 -132
rect 458 -142 463 -135
rect 568 -142 573 -113
rect 724 -118 725 -110
rect 731 -118 788 -110
rect 724 -119 732 -118
rect 458 -147 573 -142
rect 313 -156 336 -152
rect 332 -159 336 -156
rect 332 -163 488 -159
rect 251 -206 252 -200
rect 251 -207 258 -206
rect 212 -264 221 -262
rect 212 -270 271 -264
rect 201 -300 211 -295
rect 206 -340 211 -300
rect 205 -341 212 -340
rect 205 -346 206 -341
rect 211 -346 212 -341
rect 205 -347 212 -346
rect 216 -413 221 -270
rect 282 -270 316 -264
rect 332 -350 336 -163
rect 372 -183 436 -177
rect 372 -185 384 -183
rect 429 -184 445 -183
rect 371 -186 379 -185
rect 371 -192 372 -186
rect 378 -192 379 -186
rect 429 -189 449 -184
rect 484 -189 488 -163
rect 790 -173 797 -172
rect 790 -178 791 -173
rect 796 -178 797 -173
rect 790 -179 797 -178
rect 371 -193 379 -192
rect 444 -194 477 -189
rect 472 -200 477 -194
rect 483 -190 490 -189
rect 483 -195 484 -190
rect 489 -195 490 -190
rect 483 -196 490 -195
rect 518 -200 522 -188
rect 472 -204 522 -200
rect 313 -354 336 -350
rect 427 -212 487 -208
rect 313 -393 336 -392
rect 427 -393 431 -212
rect 483 -250 487 -212
rect 792 -211 795 -179
rect 792 -214 860 -211
rect 482 -251 489 -250
rect 482 -256 483 -251
rect 488 -256 489 -251
rect 482 -257 489 -256
rect 481 -311 488 -310
rect 481 -316 482 -311
rect 487 -316 488 -311
rect 481 -317 488 -316
rect 482 -333 486 -317
rect 482 -337 489 -333
rect 313 -396 431 -393
rect 332 -397 431 -396
rect 158 -414 221 -413
rect 158 -419 159 -414
rect 164 -418 221 -414
rect 164 -419 165 -418
rect 158 -420 165 -419
rect 158 -469 165 -468
rect 158 -474 159 -469
rect 164 -474 165 -469
rect 158 -475 165 -474
rect 159 -502 164 -475
rect 244 -484 251 -483
rect 234 -485 245 -484
rect 212 -489 245 -485
rect 250 -489 251 -484
rect 212 -502 218 -489
rect 244 -490 251 -489
rect 159 -507 218 -502
rect 171 -532 178 -531
rect 171 -537 172 -532
rect 177 -537 178 -532
rect 171 -538 178 -537
rect 172 -1052 177 -538
rect 212 -567 218 -507
rect 293 -567 300 -566
rect 212 -572 294 -567
rect 299 -572 300 -567
rect 212 -573 300 -572
rect 212 -695 218 -573
rect 223 -582 230 -581
rect 262 -582 269 -581
rect 223 -587 224 -582
rect 229 -587 263 -582
rect 268 -587 269 -582
rect 223 -588 230 -587
rect 252 -630 256 -587
rect 262 -588 269 -587
rect 332 -583 336 -397
rect 485 -581 489 -337
rect 313 -587 336 -583
rect 251 -637 252 -631
rect 251 -638 258 -637
rect 212 -701 271 -695
rect 332 -781 336 -587
rect 400 -585 489 -581
rect 313 -785 336 -781
rect 378 -756 385 -755
rect 378 -761 379 -756
rect 384 -761 385 -756
rect 378 -762 385 -761
rect 378 -802 384 -762
rect 212 -808 384 -802
rect 212 -916 218 -808
rect 313 -825 336 -823
rect 400 -825 404 -585
rect 313 -827 404 -825
rect 332 -829 404 -827
rect 244 -915 251 -914
rect 234 -916 245 -915
rect 212 -920 245 -916
rect 250 -920 251 -915
rect 212 -1052 218 -920
rect 244 -921 251 -920
rect 223 -1013 230 -1012
rect 262 -1013 269 -1012
rect 223 -1018 224 -1013
rect 229 -1018 263 -1013
rect 268 -1018 269 -1013
rect 223 -1019 230 -1018
rect 172 -1057 218 -1052
rect 212 -1126 218 -1057
rect 252 -1061 256 -1018
rect 262 -1019 269 -1018
rect 332 -1014 336 -829
rect 313 -1018 336 -1014
rect 251 -1068 252 -1062
rect 251 -1069 258 -1068
rect 212 -1132 271 -1126
rect 332 -1212 336 -1018
rect 313 -1216 336 -1212
<< labels >>
rlabel metal1 5 17 12 21 1 pre_A0
rlabel metal1 5 -43 12 -39 1 pre_A1
rlabel metal1 5 -103 12 -99 1 pre_A2
rlabel metal1 5 -163 12 -159 1 pre_A3
rlabel metal1 5 -223 12 -219 1 pre_A4
rlabel metal1 5 -293 12 -289 1 pre_B0
rlabel metal1 5 -353 12 -349 1 pre_B1
rlabel metal1 5 -413 12 -409 1 pre_B2
rlabel metal1 5 -473 12 -469 1 pre_B3
rlabel metal1 5 -533 12 -529 1 pre_B4
rlabel metal1 137 -534 150 -530 1 B4
rlabel metal1 137 -474 150 -470 1 B3
rlabel metal1 137 -354 150 -350 1 B1
rlabel metal1 137 -294 150 -290 1 B0
rlabel metal1 137 13 141 28 1 A0
rlabel metal1 -8 -509 -4 45 3 vdd
rlabel metal2 -1 -55 3 0 1 gnd
rlabel metal1 137 16 150 20 1 A0
rlabel metal1 137 -44 150 -40 1 A1
rlabel metal1 137 -104 150 -100 1 A2
rlabel metal1 137 -167 141 -152 1 A3
rlabel metal1 137 -227 141 -212 1 A4
rlabel metal1 137 -297 141 -282 1 B0
rlabel metal1 137 -357 141 -342 1 B1
rlabel metal1 137 -417 141 -402 1 B2
rlabel metal1 137 -477 141 -462 1 B3
rlabel metal1 137 -537 141 -522 1 B4
rlabel metal2 147 0 190 5 1 gnd
rlabel metal1 -8 41 190 45 1 vdd
rlabel metal2 339 537 346 864 1 P0
rlabel metal2 339 106 346 433 1 P1
rlabel metal2 339 -325 346 2 1 P2
rlabel metal2 339 -650 362 -643 1 P3
rlabel metal2 339 -1187 346 -860 1 P4
<< end >>
