magic
tech scmos
timestamp 1763829940
<< nwell >>
rect 49 -7 76 18
rect 49 -117 76 -92
rect 129 -112 156 -87
rect 47 -212 76 -192
rect 47 -217 74 -212
rect 127 -219 156 -197
rect 130 -222 156 -219
rect 49 -327 76 -302
<< ntransistor >>
rect 61 -28 63 -20
rect 61 -138 63 -130
rect 141 -133 143 -125
rect 61 -238 63 -230
rect 141 -243 143 -235
rect 61 -348 63 -340
<< ptransistor >>
rect 61 4 63 12
rect 61 -106 63 -98
rect 141 -101 143 -93
rect 61 -206 63 -198
rect 141 -211 143 -203
rect 61 -316 63 -308
<< ndiffusion >>
rect 60 -28 61 -20
rect 63 -28 64 -20
rect 60 -138 61 -130
rect 63 -138 64 -130
rect 140 -133 141 -125
rect 143 -133 144 -125
rect 60 -238 61 -230
rect 63 -238 64 -230
rect 140 -243 141 -235
rect 143 -243 144 -235
rect 60 -348 61 -340
rect 63 -348 64 -340
<< pdiffusion >>
rect 60 4 61 12
rect 63 4 64 12
rect 60 -106 61 -98
rect 63 -106 64 -98
rect 140 -101 141 -93
rect 143 -101 144 -93
rect 60 -206 61 -198
rect 63 -206 64 -198
rect 140 -211 141 -203
rect 143 -211 144 -203
rect 60 -316 61 -308
rect 63 -316 64 -308
<< ndcontact >>
rect 56 -28 60 -20
rect 64 -28 68 -20
rect 56 -138 60 -130
rect 64 -138 68 -130
rect 136 -133 140 -125
rect 144 -133 148 -125
rect 56 -238 60 -230
rect 64 -238 68 -230
rect 136 -243 140 -235
rect 144 -243 148 -235
rect 56 -348 60 -340
rect 64 -348 68 -340
<< pdcontact >>
rect 56 4 60 12
rect 64 4 68 12
rect 56 -106 60 -98
rect 64 -106 68 -98
rect 136 -101 140 -93
rect 144 -101 148 -93
rect 56 -206 60 -198
rect 64 -206 68 -198
rect 136 -211 140 -203
rect 144 -211 148 -203
rect 56 -316 60 -308
rect 64 -316 68 -308
<< nsubstratencontact >>
rect 68 -4 72 0
rect 148 -109 152 -105
rect 68 -114 72 -110
rect 67 -214 71 -210
rect 148 -219 152 -215
rect 68 -324 72 -320
<< polysilicon >>
rect 61 12 63 19
rect 61 -2 63 4
rect 61 -20 63 -14
rect 61 -31 63 -28
rect 61 -98 63 -90
rect 141 -93 143 -86
rect 61 -112 63 -106
rect 141 -107 143 -101
rect 61 -130 63 -124
rect 141 -125 143 -119
rect 141 -137 143 -133
rect 61 -142 63 -138
rect 61 -198 63 -191
rect 141 -203 143 -196
rect 61 -212 63 -206
rect 141 -217 143 -211
rect 61 -230 63 -224
rect 141 -235 143 -229
rect 61 -242 63 -238
rect 141 -247 143 -243
rect 61 -308 63 -301
rect 61 -322 63 -316
rect 61 -340 63 -334
rect 61 -352 63 -348
<< polycontact >>
rect 60 19 64 23
rect 60 -35 64 -31
rect 140 -86 144 -82
rect 60 -90 64 -86
rect 140 -141 144 -137
rect 60 -146 64 -142
rect 60 -191 64 -187
rect 140 -196 144 -192
rect 60 -246 64 -242
rect 140 -251 144 -247
rect 60 -301 64 -297
rect 60 -356 64 -352
<< metal1 >>
rect 60 23 64 31
rect 42 4 56 12
rect 68 4 82 12
rect 42 -20 49 4
rect 68 -11 72 -4
rect 75 -6 82 4
rect 75 -20 82 -13
rect 42 -28 56 -20
rect 68 -28 82 -20
rect 42 -60 49 -28
rect 25 -67 49 -60
rect 42 -98 49 -67
rect 60 -86 64 -35
rect 140 -82 144 -74
rect 122 -98 136 -93
rect 42 -106 56 -98
rect 68 -101 136 -98
rect 148 -101 162 -93
rect 68 -106 129 -101
rect 42 -130 49 -106
rect 68 -121 72 -114
rect 75 -130 82 -106
rect 42 -138 56 -130
rect 68 -138 82 -130
rect 122 -125 129 -106
rect 148 -116 152 -109
rect 155 -125 162 -101
rect 122 -133 136 -125
rect 148 -133 162 -125
rect 60 -187 64 -146
rect 75 -192 82 -138
rect 74 -198 82 -192
rect 140 -192 144 -141
rect 155 -164 162 -133
rect 155 -171 179 -164
rect 42 -206 56 -198
rect 68 -206 82 -198
rect 155 -203 162 -171
rect 42 -230 49 -206
rect 67 -221 71 -214
rect 74 -217 82 -206
rect 75 -230 82 -217
rect 42 -238 56 -230
rect 68 -238 82 -230
rect 122 -211 136 -203
rect 148 -211 162 -203
rect 122 -220 129 -211
rect 148 -226 152 -219
rect 122 -235 129 -227
rect 155 -235 162 -211
rect 42 -271 49 -238
rect 25 -278 49 -271
rect 42 -308 49 -278
rect 122 -243 136 -235
rect 148 -243 162 -235
rect 60 -297 64 -246
rect 140 -257 144 -251
rect 42 -316 56 -308
rect 68 -316 82 -308
rect 42 -340 49 -316
rect 68 -331 72 -324
rect 75 -326 82 -316
rect 75 -340 82 -333
rect 42 -348 56 -340
rect 68 -348 82 -340
rect 60 -362 64 -356
<< m2contact >>
rect 75 -13 82 -6
rect 122 -227 129 -220
rect 75 -333 82 -326
<< metal2 >>
rect 82 -13 99 -6
rect 92 -220 99 -13
rect 92 -227 122 -220
rect 92 -326 99 -227
rect 82 -333 99 -326
<< labels >>
rlabel metal1 25 -278 49 -271 1 B
rlabel metal1 155 -171 179 -164 1 out_XOR_3
rlabel metal1 68 -11 72 0 1 vdd
rlabel metal1 68 -121 72 -110 1 vdd
rlabel metal1 67 -221 71 -210 1 vdd
rlabel metal1 68 -331 72 -320 1 vdd
rlabel metal1 148 -226 152 -215 1 vdd
rlabel metal1 148 -116 152 -105 1 vdd
rlabel metal1 25 -67 49 -60 1 B_bar
rlabel metal1 42 -348 49 -198 1 B
rlabel metal1 60 19 64 31 1 A
rlabel metal1 60 -90 64 -31 1 A_bar
rlabel metal1 60 -191 64 -142 1 A
rlabel metal1 60 -301 64 -242 1 A_bar
rlabel metal1 60 -362 64 -352 1 A
rlabel metal1 140 -257 144 -247 1 C
rlabel metal1 140 -196 144 -137 1 C_bar
rlabel metal1 140 -86 144 -74 1 C
<< end >>
