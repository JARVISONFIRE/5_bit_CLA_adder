magic
tech scmos
timestamp 1764731542
<< nwell >>
rect 239 807 266 832
rect 185 753 210 776
rect 239 697 266 722
rect 195 605 220 628
rect 237 602 266 622
rect 237 597 264 602
rect 239 487 266 512
rect 239 395 266 420
rect 185 341 210 364
rect 239 285 266 310
rect 195 193 220 216
rect 237 190 266 210
rect 237 185 264 190
rect 239 75 266 100
rect 3 20 35 40
rect 46 20 70 40
rect 84 20 108 40
rect 122 21 147 44
rect 3 -34 35 -14
rect 46 -34 70 -14
rect 84 -34 108 -14
rect 122 -33 147 -10
rect 240 -13 267 12
rect 3 -88 35 -68
rect 46 -88 70 -68
rect 84 -88 108 -68
rect 122 -87 147 -64
rect 186 -67 211 -44
rect 371 -59 403 -39
rect 413 -58 438 -35
rect 3 -142 35 -122
rect 46 -142 70 -122
rect 84 -142 108 -122
rect 122 -141 147 -118
rect 240 -123 267 -98
rect 371 -110 403 -90
rect 413 -109 438 -86
rect 371 -161 403 -141
rect 413 -160 438 -137
rect 3 -196 35 -176
rect 46 -196 70 -176
rect 84 -196 108 -176
rect 122 -195 147 -172
rect 196 -215 221 -192
rect 238 -218 267 -198
rect 371 -212 403 -192
rect 413 -211 438 -188
rect 238 -223 265 -218
rect 4 -266 36 -246
rect 47 -266 71 -246
rect 85 -266 109 -246
rect 123 -265 148 -242
rect 371 -263 403 -243
rect 413 -262 438 -239
rect 4 -320 36 -300
rect 47 -320 71 -300
rect 85 -320 109 -300
rect 123 -319 148 -296
rect 240 -333 267 -308
rect 4 -374 36 -354
rect 47 -374 71 -354
rect 85 -374 109 -354
rect 123 -373 148 -350
rect 4 -428 36 -408
rect 47 -428 71 -408
rect 85 -428 109 -408
rect 123 -427 148 -404
rect 240 -416 267 -391
rect 4 -482 36 -462
rect 47 -482 71 -462
rect 85 -482 109 -462
rect 123 -481 148 -458
rect 186 -470 211 -447
rect 240 -526 267 -501
rect 196 -618 221 -595
rect 238 -621 267 -601
rect 238 -626 265 -621
rect 240 -736 267 -711
rect 240 -821 267 -796
rect 186 -875 211 -852
rect 240 -931 267 -906
rect 196 -1023 221 -1000
rect 238 -1026 267 -1006
rect 238 -1031 265 -1026
rect 240 -1141 267 -1116
<< ntransistor >>
rect 251 786 253 794
rect 197 741 199 745
rect 251 676 253 684
rect 207 593 209 597
rect 251 576 253 584
rect 251 466 253 474
rect 251 374 253 382
rect 197 329 199 333
rect 251 264 253 272
rect 207 181 209 185
rect 251 164 253 172
rect 251 54 253 62
rect 14 9 16 13
rect 57 9 59 13
rect 65 9 67 13
rect 95 9 97 13
rect 103 9 105 13
rect 134 9 136 13
rect 252 -34 254 -26
rect 14 -45 16 -41
rect 57 -45 59 -41
rect 65 -45 67 -41
rect 95 -45 97 -41
rect 103 -45 105 -41
rect 134 -45 136 -41
rect 382 -70 384 -66
rect 390 -70 392 -66
rect 425 -70 427 -66
rect 198 -79 200 -75
rect 14 -99 16 -95
rect 57 -99 59 -95
rect 65 -99 67 -95
rect 95 -99 97 -95
rect 103 -99 105 -95
rect 134 -99 136 -95
rect 382 -121 384 -117
rect 390 -121 392 -117
rect 425 -121 427 -117
rect 252 -144 254 -136
rect 14 -153 16 -149
rect 57 -153 59 -149
rect 65 -153 67 -149
rect 95 -153 97 -149
rect 103 -153 105 -149
rect 134 -153 136 -149
rect 382 -172 384 -168
rect 390 -172 392 -168
rect 425 -172 427 -168
rect 14 -207 16 -203
rect 57 -207 59 -203
rect 65 -207 67 -203
rect 95 -207 97 -203
rect 103 -207 105 -203
rect 134 -207 136 -203
rect 382 -223 384 -219
rect 390 -223 392 -219
rect 425 -223 427 -219
rect 208 -227 210 -223
rect 252 -244 254 -236
rect 15 -277 17 -273
rect 58 -277 60 -273
rect 66 -277 68 -273
rect 96 -277 98 -273
rect 104 -277 106 -273
rect 135 -277 137 -273
rect 382 -274 384 -270
rect 390 -274 392 -270
rect 425 -274 427 -270
rect 15 -331 17 -327
rect 58 -331 60 -327
rect 66 -331 68 -327
rect 96 -331 98 -327
rect 104 -331 106 -327
rect 135 -331 137 -327
rect 252 -354 254 -346
rect 15 -385 17 -381
rect 58 -385 60 -381
rect 66 -385 68 -381
rect 96 -385 98 -381
rect 104 -385 106 -381
rect 135 -385 137 -381
rect 15 -439 17 -435
rect 58 -439 60 -435
rect 66 -439 68 -435
rect 96 -439 98 -435
rect 104 -439 106 -435
rect 135 -439 137 -435
rect 252 -437 254 -429
rect 198 -482 200 -478
rect 15 -493 17 -489
rect 58 -493 60 -489
rect 66 -493 68 -489
rect 96 -493 98 -489
rect 104 -493 106 -489
rect 135 -493 137 -489
rect 252 -547 254 -539
rect 208 -630 210 -626
rect 252 -647 254 -639
rect 252 -757 254 -749
rect 252 -842 254 -834
rect 198 -887 200 -883
rect 252 -952 254 -944
rect 208 -1035 210 -1031
rect 252 -1052 254 -1044
rect 252 -1162 254 -1154
<< ptransistor >>
rect 251 818 253 826
rect 197 760 199 768
rect 251 708 253 716
rect 207 612 209 620
rect 251 608 253 616
rect 251 498 253 506
rect 251 406 253 414
rect 197 348 199 356
rect 251 296 253 304
rect 207 200 209 208
rect 251 196 253 204
rect 251 86 253 94
rect 14 26 16 34
rect 22 26 24 34
rect 57 26 59 34
rect 95 26 97 34
rect 134 28 136 36
rect 252 -2 254 6
rect 14 -28 16 -20
rect 22 -28 24 -20
rect 57 -28 59 -20
rect 95 -28 97 -20
rect 134 -26 136 -18
rect 198 -60 200 -52
rect 382 -53 384 -45
rect 390 -53 392 -45
rect 425 -51 427 -43
rect 14 -82 16 -74
rect 22 -82 24 -74
rect 57 -82 59 -74
rect 95 -82 97 -74
rect 134 -80 136 -72
rect 382 -104 384 -96
rect 390 -104 392 -96
rect 425 -102 427 -94
rect 252 -112 254 -104
rect 14 -136 16 -128
rect 22 -136 24 -128
rect 57 -136 59 -128
rect 95 -136 97 -128
rect 134 -134 136 -126
rect 382 -155 384 -147
rect 390 -155 392 -147
rect 425 -153 427 -145
rect 14 -190 16 -182
rect 22 -190 24 -182
rect 57 -190 59 -182
rect 95 -190 97 -182
rect 134 -188 136 -180
rect 208 -208 210 -200
rect 252 -212 254 -204
rect 382 -206 384 -198
rect 390 -206 392 -198
rect 425 -204 427 -196
rect 15 -260 17 -252
rect 23 -260 25 -252
rect 58 -260 60 -252
rect 96 -260 98 -252
rect 135 -258 137 -250
rect 382 -257 384 -249
rect 390 -257 392 -249
rect 425 -255 427 -247
rect 15 -314 17 -306
rect 23 -314 25 -306
rect 58 -314 60 -306
rect 96 -314 98 -306
rect 135 -312 137 -304
rect 252 -322 254 -314
rect 15 -368 17 -360
rect 23 -368 25 -360
rect 58 -368 60 -360
rect 96 -368 98 -360
rect 135 -366 137 -358
rect 252 -405 254 -397
rect 15 -422 17 -414
rect 23 -422 25 -414
rect 58 -422 60 -414
rect 96 -422 98 -414
rect 135 -420 137 -412
rect 198 -463 200 -455
rect 15 -476 17 -468
rect 23 -476 25 -468
rect 58 -476 60 -468
rect 96 -476 98 -468
rect 135 -474 137 -466
rect 252 -515 254 -507
rect 208 -611 210 -603
rect 252 -615 254 -607
rect 252 -725 254 -717
rect 252 -810 254 -802
rect 198 -868 200 -860
rect 252 -920 254 -912
rect 208 -1016 210 -1008
rect 252 -1020 254 -1012
rect 252 -1130 254 -1122
<< ndiffusion >>
rect 250 786 251 794
rect 253 786 254 794
rect 196 741 197 745
rect 199 741 200 745
rect 250 676 251 684
rect 253 676 254 684
rect 206 593 207 597
rect 209 593 210 597
rect 250 576 251 584
rect 253 576 254 584
rect 250 466 251 474
rect 253 466 254 474
rect 250 374 251 382
rect 253 374 254 382
rect 196 329 197 333
rect 199 329 200 333
rect 250 264 251 272
rect 253 264 254 272
rect 206 181 207 185
rect 209 181 210 185
rect 250 164 251 172
rect 253 164 254 172
rect 250 54 251 62
rect 253 54 254 62
rect 13 9 14 13
rect 16 9 17 13
rect 56 9 57 13
rect 59 9 60 13
rect 64 9 65 13
rect 67 9 68 13
rect 94 9 95 13
rect 97 9 98 13
rect 102 9 103 13
rect 105 9 106 13
rect 133 9 134 13
rect 136 9 137 13
rect 251 -34 252 -26
rect 254 -34 255 -26
rect 13 -45 14 -41
rect 16 -45 17 -41
rect 56 -45 57 -41
rect 59 -45 60 -41
rect 64 -45 65 -41
rect 67 -45 68 -41
rect 94 -45 95 -41
rect 97 -45 98 -41
rect 102 -45 103 -41
rect 105 -45 106 -41
rect 133 -45 134 -41
rect 136 -45 137 -41
rect 381 -70 382 -66
rect 384 -70 385 -66
rect 389 -70 390 -66
rect 392 -70 393 -66
rect 424 -70 425 -66
rect 427 -70 428 -66
rect 197 -79 198 -75
rect 200 -79 201 -75
rect 13 -99 14 -95
rect 16 -99 17 -95
rect 56 -99 57 -95
rect 59 -99 60 -95
rect 64 -99 65 -95
rect 67 -99 68 -95
rect 94 -99 95 -95
rect 97 -99 98 -95
rect 102 -99 103 -95
rect 105 -99 106 -95
rect 133 -99 134 -95
rect 136 -99 137 -95
rect 381 -121 382 -117
rect 384 -121 385 -117
rect 389 -121 390 -117
rect 392 -121 393 -117
rect 424 -121 425 -117
rect 427 -121 428 -117
rect 251 -144 252 -136
rect 254 -144 255 -136
rect 13 -153 14 -149
rect 16 -153 17 -149
rect 56 -153 57 -149
rect 59 -153 60 -149
rect 64 -153 65 -149
rect 67 -153 68 -149
rect 94 -153 95 -149
rect 97 -153 98 -149
rect 102 -153 103 -149
rect 105 -153 106 -149
rect 133 -153 134 -149
rect 136 -153 137 -149
rect 381 -172 382 -168
rect 384 -172 385 -168
rect 389 -172 390 -168
rect 392 -172 393 -168
rect 424 -172 425 -168
rect 427 -172 428 -168
rect 13 -207 14 -203
rect 16 -207 17 -203
rect 56 -207 57 -203
rect 59 -207 60 -203
rect 64 -207 65 -203
rect 67 -207 68 -203
rect 94 -207 95 -203
rect 97 -207 98 -203
rect 102 -207 103 -203
rect 105 -207 106 -203
rect 133 -207 134 -203
rect 136 -207 137 -203
rect 381 -223 382 -219
rect 384 -223 385 -219
rect 389 -223 390 -219
rect 392 -223 393 -219
rect 424 -223 425 -219
rect 427 -223 428 -219
rect 207 -227 208 -223
rect 210 -227 211 -223
rect 251 -244 252 -236
rect 254 -244 255 -236
rect 14 -277 15 -273
rect 17 -277 18 -273
rect 57 -277 58 -273
rect 60 -277 61 -273
rect 65 -277 66 -273
rect 68 -277 69 -273
rect 95 -277 96 -273
rect 98 -277 99 -273
rect 103 -277 104 -273
rect 106 -277 107 -273
rect 134 -277 135 -273
rect 137 -277 138 -273
rect 381 -274 382 -270
rect 384 -274 385 -270
rect 389 -274 390 -270
rect 392 -274 393 -270
rect 424 -274 425 -270
rect 427 -274 428 -270
rect 14 -331 15 -327
rect 17 -331 18 -327
rect 57 -331 58 -327
rect 60 -331 61 -327
rect 65 -331 66 -327
rect 68 -331 69 -327
rect 95 -331 96 -327
rect 98 -331 99 -327
rect 103 -331 104 -327
rect 106 -331 107 -327
rect 134 -331 135 -327
rect 137 -331 138 -327
rect 251 -354 252 -346
rect 254 -354 255 -346
rect 14 -385 15 -381
rect 17 -385 18 -381
rect 57 -385 58 -381
rect 60 -385 61 -381
rect 65 -385 66 -381
rect 68 -385 69 -381
rect 95 -385 96 -381
rect 98 -385 99 -381
rect 103 -385 104 -381
rect 106 -385 107 -381
rect 134 -385 135 -381
rect 137 -385 138 -381
rect 14 -439 15 -435
rect 17 -439 18 -435
rect 57 -439 58 -435
rect 60 -439 61 -435
rect 65 -439 66 -435
rect 68 -439 69 -435
rect 95 -439 96 -435
rect 98 -439 99 -435
rect 103 -439 104 -435
rect 106 -439 107 -435
rect 134 -439 135 -435
rect 137 -439 138 -435
rect 251 -437 252 -429
rect 254 -437 255 -429
rect 197 -482 198 -478
rect 200 -482 201 -478
rect 14 -493 15 -489
rect 17 -493 18 -489
rect 57 -493 58 -489
rect 60 -493 61 -489
rect 65 -493 66 -489
rect 68 -493 69 -489
rect 95 -493 96 -489
rect 98 -493 99 -489
rect 103 -493 104 -489
rect 106 -493 107 -489
rect 134 -493 135 -489
rect 137 -493 138 -489
rect 251 -547 252 -539
rect 254 -547 255 -539
rect 207 -630 208 -626
rect 210 -630 211 -626
rect 251 -647 252 -639
rect 254 -647 255 -639
rect 251 -757 252 -749
rect 254 -757 255 -749
rect 251 -842 252 -834
rect 254 -842 255 -834
rect 197 -887 198 -883
rect 200 -887 201 -883
rect 251 -952 252 -944
rect 254 -952 255 -944
rect 207 -1035 208 -1031
rect 210 -1035 211 -1031
rect 251 -1052 252 -1044
rect 254 -1052 255 -1044
rect 251 -1162 252 -1154
rect 254 -1162 255 -1154
<< pdiffusion >>
rect 250 818 251 826
rect 253 818 254 826
rect 196 760 197 768
rect 199 760 200 768
rect 250 708 251 716
rect 253 708 254 716
rect 206 612 207 620
rect 209 612 210 620
rect 250 608 251 616
rect 253 608 254 616
rect 250 498 251 506
rect 253 498 254 506
rect 250 406 251 414
rect 253 406 254 414
rect 196 348 197 356
rect 199 348 200 356
rect 250 296 251 304
rect 253 296 254 304
rect 206 200 207 208
rect 209 200 210 208
rect 250 196 251 204
rect 253 196 254 204
rect 250 86 251 94
rect 253 86 254 94
rect 13 26 14 34
rect 16 26 17 34
rect 21 26 22 34
rect 24 26 25 34
rect 56 26 57 34
rect 59 26 60 34
rect 94 26 95 34
rect 97 26 98 34
rect 133 28 134 36
rect 136 28 137 36
rect 251 -2 252 6
rect 254 -2 255 6
rect 13 -28 14 -20
rect 16 -28 17 -20
rect 21 -28 22 -20
rect 24 -28 25 -20
rect 56 -28 57 -20
rect 59 -28 60 -20
rect 94 -28 95 -20
rect 97 -28 98 -20
rect 133 -26 134 -18
rect 136 -26 137 -18
rect 197 -60 198 -52
rect 200 -60 201 -52
rect 381 -53 382 -45
rect 384 -53 385 -45
rect 389 -53 390 -45
rect 392 -53 393 -45
rect 424 -51 425 -43
rect 427 -51 428 -43
rect 13 -82 14 -74
rect 16 -82 17 -74
rect 21 -82 22 -74
rect 24 -82 25 -74
rect 56 -82 57 -74
rect 59 -82 60 -74
rect 94 -82 95 -74
rect 97 -82 98 -74
rect 133 -80 134 -72
rect 136 -80 137 -72
rect 381 -104 382 -96
rect 384 -104 385 -96
rect 389 -104 390 -96
rect 392 -104 393 -96
rect 424 -102 425 -94
rect 427 -102 428 -94
rect 251 -112 252 -104
rect 254 -112 255 -104
rect 13 -136 14 -128
rect 16 -136 17 -128
rect 21 -136 22 -128
rect 24 -136 25 -128
rect 56 -136 57 -128
rect 59 -136 60 -128
rect 94 -136 95 -128
rect 97 -136 98 -128
rect 133 -134 134 -126
rect 136 -134 137 -126
rect 381 -155 382 -147
rect 384 -155 385 -147
rect 389 -155 390 -147
rect 392 -155 393 -147
rect 424 -153 425 -145
rect 427 -153 428 -145
rect 13 -190 14 -182
rect 16 -190 17 -182
rect 21 -190 22 -182
rect 24 -190 25 -182
rect 56 -190 57 -182
rect 59 -190 60 -182
rect 94 -190 95 -182
rect 97 -190 98 -182
rect 133 -188 134 -180
rect 136 -188 137 -180
rect 207 -208 208 -200
rect 210 -208 211 -200
rect 251 -212 252 -204
rect 254 -212 255 -204
rect 381 -206 382 -198
rect 384 -206 385 -198
rect 389 -206 390 -198
rect 392 -206 393 -198
rect 424 -204 425 -196
rect 427 -204 428 -196
rect 14 -260 15 -252
rect 17 -260 18 -252
rect 22 -260 23 -252
rect 25 -260 26 -252
rect 57 -260 58 -252
rect 60 -260 61 -252
rect 95 -260 96 -252
rect 98 -260 99 -252
rect 134 -258 135 -250
rect 137 -258 138 -250
rect 381 -257 382 -249
rect 384 -257 385 -249
rect 389 -257 390 -249
rect 392 -257 393 -249
rect 424 -255 425 -247
rect 427 -255 428 -247
rect 14 -314 15 -306
rect 17 -314 18 -306
rect 22 -314 23 -306
rect 25 -314 26 -306
rect 57 -314 58 -306
rect 60 -314 61 -306
rect 95 -314 96 -306
rect 98 -314 99 -306
rect 134 -312 135 -304
rect 137 -312 138 -304
rect 251 -322 252 -314
rect 254 -322 255 -314
rect 14 -368 15 -360
rect 17 -368 18 -360
rect 22 -368 23 -360
rect 25 -368 26 -360
rect 57 -368 58 -360
rect 60 -368 61 -360
rect 95 -368 96 -360
rect 98 -368 99 -360
rect 134 -366 135 -358
rect 137 -366 138 -358
rect 251 -405 252 -397
rect 254 -405 255 -397
rect 14 -422 15 -414
rect 17 -422 18 -414
rect 22 -422 23 -414
rect 25 -422 26 -414
rect 57 -422 58 -414
rect 60 -422 61 -414
rect 95 -422 96 -414
rect 98 -422 99 -414
rect 134 -420 135 -412
rect 137 -420 138 -412
rect 197 -463 198 -455
rect 200 -463 201 -455
rect 14 -476 15 -468
rect 17 -476 18 -468
rect 22 -476 23 -468
rect 25 -476 26 -468
rect 57 -476 58 -468
rect 60 -476 61 -468
rect 95 -476 96 -468
rect 98 -476 99 -468
rect 134 -474 135 -466
rect 137 -474 138 -466
rect 251 -515 252 -507
rect 254 -515 255 -507
rect 207 -611 208 -603
rect 210 -611 211 -603
rect 251 -615 252 -607
rect 254 -615 255 -607
rect 251 -725 252 -717
rect 254 -725 255 -717
rect 251 -810 252 -802
rect 254 -810 255 -802
rect 197 -868 198 -860
rect 200 -868 201 -860
rect 251 -920 252 -912
rect 254 -920 255 -912
rect 207 -1016 208 -1008
rect 210 -1016 211 -1008
rect 251 -1020 252 -1012
rect 254 -1020 255 -1012
rect 251 -1130 252 -1122
rect 254 -1130 255 -1122
<< ndcontact >>
rect 246 786 250 794
rect 254 786 258 794
rect 192 741 196 745
rect 200 741 204 745
rect 246 676 250 684
rect 254 676 258 684
rect 202 593 206 597
rect 210 593 214 597
rect 246 576 250 584
rect 254 576 258 584
rect 246 466 250 474
rect 254 466 258 474
rect 246 374 250 382
rect 254 374 258 382
rect 192 329 196 333
rect 200 329 204 333
rect 246 264 250 272
rect 254 264 258 272
rect 202 181 206 185
rect 210 181 214 185
rect 246 164 250 172
rect 254 164 258 172
rect 246 54 250 62
rect 254 54 258 62
rect 9 9 13 13
rect 17 9 21 13
rect 52 9 56 13
rect 60 9 64 13
rect 68 9 72 13
rect 90 9 94 13
rect 98 9 102 13
rect 106 9 110 13
rect 129 9 133 13
rect 137 9 141 13
rect 247 -34 251 -26
rect 255 -34 259 -26
rect 9 -45 13 -41
rect 17 -45 21 -41
rect 52 -45 56 -41
rect 60 -45 64 -41
rect 68 -45 72 -41
rect 90 -45 94 -41
rect 98 -45 102 -41
rect 106 -45 110 -41
rect 129 -45 133 -41
rect 137 -45 141 -41
rect 377 -70 381 -66
rect 385 -70 389 -66
rect 393 -70 397 -66
rect 420 -70 424 -66
rect 428 -70 432 -66
rect 193 -79 197 -75
rect 201 -79 205 -75
rect 9 -99 13 -95
rect 17 -99 21 -95
rect 52 -99 56 -95
rect 60 -99 64 -95
rect 68 -99 72 -95
rect 90 -99 94 -95
rect 98 -99 102 -95
rect 106 -99 110 -95
rect 129 -99 133 -95
rect 137 -99 141 -95
rect 377 -121 381 -117
rect 385 -121 389 -117
rect 393 -121 397 -117
rect 420 -121 424 -117
rect 428 -121 432 -117
rect 247 -144 251 -136
rect 255 -144 259 -136
rect 9 -153 13 -149
rect 17 -153 21 -149
rect 52 -153 56 -149
rect 60 -153 64 -149
rect 68 -153 72 -149
rect 90 -153 94 -149
rect 98 -153 102 -149
rect 106 -153 110 -149
rect 129 -153 133 -149
rect 137 -153 141 -149
rect 377 -172 381 -168
rect 385 -172 389 -168
rect 393 -172 397 -168
rect 420 -172 424 -168
rect 428 -172 432 -168
rect 9 -207 13 -203
rect 17 -207 21 -203
rect 52 -207 56 -203
rect 60 -207 64 -203
rect 68 -207 72 -203
rect 90 -207 94 -203
rect 98 -207 102 -203
rect 106 -207 110 -203
rect 129 -207 133 -203
rect 137 -207 141 -203
rect 377 -223 381 -219
rect 385 -223 389 -219
rect 393 -223 397 -219
rect 420 -223 424 -219
rect 428 -223 432 -219
rect 203 -227 207 -223
rect 211 -227 215 -223
rect 247 -244 251 -236
rect 255 -244 259 -236
rect 10 -277 14 -273
rect 18 -277 22 -273
rect 53 -277 57 -273
rect 61 -277 65 -273
rect 69 -277 73 -273
rect 91 -277 95 -273
rect 99 -277 103 -273
rect 107 -277 111 -273
rect 130 -277 134 -273
rect 138 -277 142 -273
rect 377 -274 381 -270
rect 385 -274 389 -270
rect 393 -274 397 -270
rect 420 -274 424 -270
rect 428 -274 432 -270
rect 10 -331 14 -327
rect 18 -331 22 -327
rect 53 -331 57 -327
rect 61 -331 65 -327
rect 69 -331 73 -327
rect 91 -331 95 -327
rect 99 -331 103 -327
rect 107 -331 111 -327
rect 130 -331 134 -327
rect 138 -331 142 -327
rect 247 -354 251 -346
rect 255 -354 259 -346
rect 10 -385 14 -381
rect 18 -385 22 -381
rect 53 -385 57 -381
rect 61 -385 65 -381
rect 69 -385 73 -381
rect 91 -385 95 -381
rect 99 -385 103 -381
rect 107 -385 111 -381
rect 130 -385 134 -381
rect 138 -385 142 -381
rect 10 -439 14 -435
rect 18 -439 22 -435
rect 53 -439 57 -435
rect 61 -439 65 -435
rect 69 -439 73 -435
rect 91 -439 95 -435
rect 99 -439 103 -435
rect 107 -439 111 -435
rect 130 -439 134 -435
rect 138 -439 142 -435
rect 247 -437 251 -429
rect 255 -437 259 -429
rect 193 -482 197 -478
rect 201 -482 205 -478
rect 10 -493 14 -489
rect 18 -493 22 -489
rect 53 -493 57 -489
rect 61 -493 65 -489
rect 69 -493 73 -489
rect 91 -493 95 -489
rect 99 -493 103 -489
rect 107 -493 111 -489
rect 130 -493 134 -489
rect 138 -493 142 -489
rect 247 -547 251 -539
rect 255 -547 259 -539
rect 203 -630 207 -626
rect 211 -630 215 -626
rect 247 -647 251 -639
rect 255 -647 259 -639
rect 247 -757 251 -749
rect 255 -757 259 -749
rect 247 -842 251 -834
rect 255 -842 259 -834
rect 193 -887 197 -883
rect 201 -887 205 -883
rect 247 -952 251 -944
rect 255 -952 259 -944
rect 203 -1035 207 -1031
rect 211 -1035 215 -1031
rect 247 -1052 251 -1044
rect 255 -1052 259 -1044
rect 247 -1162 251 -1154
rect 255 -1162 259 -1154
<< pdcontact >>
rect 246 818 250 826
rect 254 818 258 826
rect 192 760 196 768
rect 200 760 204 768
rect 246 708 250 716
rect 254 708 258 716
rect 202 612 206 620
rect 210 612 214 620
rect 246 608 250 616
rect 254 608 258 616
rect 246 498 250 506
rect 254 498 258 506
rect 246 406 250 414
rect 254 406 258 414
rect 192 348 196 356
rect 200 348 204 356
rect 246 296 250 304
rect 254 296 258 304
rect 202 200 206 208
rect 210 200 214 208
rect 246 196 250 204
rect 254 196 258 204
rect 246 86 250 94
rect 254 86 258 94
rect 9 26 13 34
rect 17 26 21 34
rect 25 26 29 34
rect 52 26 56 34
rect 60 26 64 34
rect 90 26 94 34
rect 98 26 102 34
rect 129 28 133 36
rect 137 28 141 36
rect 247 -2 251 6
rect 255 -2 259 6
rect 9 -28 13 -20
rect 17 -28 21 -20
rect 25 -28 29 -20
rect 52 -28 56 -20
rect 60 -28 64 -20
rect 90 -28 94 -20
rect 98 -28 102 -20
rect 129 -26 133 -18
rect 137 -26 141 -18
rect 193 -60 197 -52
rect 201 -60 205 -52
rect 377 -53 381 -45
rect 385 -53 389 -45
rect 393 -53 397 -45
rect 420 -51 424 -43
rect 428 -51 432 -43
rect 9 -82 13 -74
rect 17 -82 21 -74
rect 25 -82 29 -74
rect 52 -82 56 -74
rect 60 -82 64 -74
rect 90 -82 94 -74
rect 98 -82 102 -74
rect 129 -80 133 -72
rect 137 -80 141 -72
rect 377 -104 381 -96
rect 385 -104 389 -96
rect 393 -104 397 -96
rect 420 -102 424 -94
rect 428 -102 432 -94
rect 247 -112 251 -104
rect 255 -112 259 -104
rect 9 -136 13 -128
rect 17 -136 21 -128
rect 25 -136 29 -128
rect 52 -136 56 -128
rect 60 -136 64 -128
rect 90 -136 94 -128
rect 98 -136 102 -128
rect 129 -134 133 -126
rect 137 -134 141 -126
rect 377 -155 381 -147
rect 385 -155 389 -147
rect 393 -155 397 -147
rect 420 -153 424 -145
rect 428 -153 432 -145
rect 9 -190 13 -182
rect 17 -190 21 -182
rect 25 -190 29 -182
rect 52 -190 56 -182
rect 60 -190 64 -182
rect 90 -190 94 -182
rect 98 -190 102 -182
rect 129 -188 133 -180
rect 137 -188 141 -180
rect 203 -208 207 -200
rect 211 -208 215 -200
rect 247 -212 251 -204
rect 255 -212 259 -204
rect 377 -206 381 -198
rect 385 -206 389 -198
rect 393 -206 397 -198
rect 420 -204 424 -196
rect 428 -204 432 -196
rect 10 -260 14 -252
rect 18 -260 22 -252
rect 26 -260 30 -252
rect 53 -260 57 -252
rect 61 -260 65 -252
rect 91 -260 95 -252
rect 99 -260 103 -252
rect 130 -258 134 -250
rect 138 -258 142 -250
rect 377 -257 381 -249
rect 385 -257 389 -249
rect 393 -257 397 -249
rect 420 -255 424 -247
rect 428 -255 432 -247
rect 10 -314 14 -306
rect 18 -314 22 -306
rect 26 -314 30 -306
rect 53 -314 57 -306
rect 61 -314 65 -306
rect 91 -314 95 -306
rect 99 -314 103 -306
rect 130 -312 134 -304
rect 138 -312 142 -304
rect 247 -322 251 -314
rect 255 -322 259 -314
rect 10 -368 14 -360
rect 18 -368 22 -360
rect 26 -368 30 -360
rect 53 -368 57 -360
rect 61 -368 65 -360
rect 91 -368 95 -360
rect 99 -368 103 -360
rect 130 -366 134 -358
rect 138 -366 142 -358
rect 247 -405 251 -397
rect 255 -405 259 -397
rect 10 -422 14 -414
rect 18 -422 22 -414
rect 26 -422 30 -414
rect 53 -422 57 -414
rect 61 -422 65 -414
rect 91 -422 95 -414
rect 99 -422 103 -414
rect 130 -420 134 -412
rect 138 -420 142 -412
rect 193 -463 197 -455
rect 201 -463 205 -455
rect 10 -476 14 -468
rect 18 -476 22 -468
rect 26 -476 30 -468
rect 53 -476 57 -468
rect 61 -476 65 -468
rect 91 -476 95 -468
rect 99 -476 103 -468
rect 130 -474 134 -466
rect 138 -474 142 -466
rect 247 -515 251 -507
rect 255 -515 259 -507
rect 203 -611 207 -603
rect 211 -611 215 -603
rect 247 -615 251 -607
rect 255 -615 259 -607
rect 247 -725 251 -717
rect 255 -725 259 -717
rect 247 -810 251 -802
rect 255 -810 259 -802
rect 193 -868 197 -860
rect 201 -868 205 -860
rect 247 -920 251 -912
rect 255 -920 259 -912
rect 203 -1016 207 -1008
rect 211 -1016 215 -1008
rect 247 -1020 251 -1012
rect 255 -1020 259 -1012
rect 247 -1130 251 -1122
rect 255 -1130 259 -1122
<< nsubstratencontact >>
rect 258 810 262 814
rect 258 700 262 704
rect 257 600 261 604
rect 258 490 262 494
rect 258 398 262 402
rect 258 288 262 292
rect 257 188 261 192
rect 258 78 262 82
rect 259 -10 263 -6
rect 259 -120 263 -116
rect 258 -220 262 -216
rect 259 -330 263 -326
rect 259 -413 263 -409
rect 259 -523 263 -519
rect 258 -623 262 -619
rect 259 -733 263 -729
rect 259 -818 263 -814
rect 259 -928 263 -924
rect 258 -1028 262 -1024
rect 259 -1138 263 -1134
<< polysilicon >>
rect 251 826 253 833
rect 251 812 253 818
rect 251 794 253 800
rect 251 783 253 786
rect 197 768 199 771
rect 197 745 199 760
rect 197 738 199 741
rect 251 716 253 724
rect 251 702 253 708
rect 251 684 253 690
rect 251 672 253 676
rect 207 620 209 623
rect 251 616 253 623
rect 207 597 209 612
rect 251 602 253 608
rect 207 590 209 593
rect 251 584 253 590
rect 251 572 253 576
rect 251 506 253 513
rect 251 492 253 498
rect 251 474 253 480
rect 251 462 253 466
rect 251 414 253 421
rect 251 400 253 406
rect 251 382 253 388
rect 251 371 253 374
rect 197 356 199 359
rect 197 333 199 348
rect 197 326 199 329
rect 251 304 253 312
rect 251 290 253 296
rect 251 272 253 278
rect 251 260 253 264
rect 207 208 209 211
rect 251 204 253 211
rect 207 185 209 200
rect 251 190 253 196
rect 207 178 209 181
rect 251 172 253 178
rect 251 160 253 164
rect 251 94 253 101
rect 251 80 253 86
rect 251 62 253 68
rect 251 50 253 54
rect 14 34 16 38
rect 22 36 32 38
rect 22 34 24 36
rect 57 34 59 38
rect 95 34 97 38
rect 134 36 136 39
rect 14 21 16 26
rect 22 23 24 26
rect 57 20 59 26
rect 95 20 97 26
rect 14 13 16 17
rect 57 13 59 16
rect 65 15 75 17
rect 65 13 67 15
rect 95 13 97 16
rect 103 15 113 17
rect 103 13 105 15
rect 134 13 136 28
rect 14 5 16 9
rect 57 5 59 9
rect 65 5 67 9
rect 95 5 97 9
rect 103 5 105 9
rect 134 6 136 9
rect 252 6 254 13
rect 252 -8 254 -2
rect 14 -20 16 -16
rect 22 -18 32 -16
rect 22 -20 24 -18
rect 57 -20 59 -16
rect 95 -20 97 -16
rect 134 -18 136 -15
rect 252 -26 254 -20
rect 14 -33 16 -28
rect 22 -31 24 -28
rect 57 -34 59 -28
rect 95 -34 97 -28
rect 14 -41 16 -37
rect 57 -41 59 -38
rect 65 -39 75 -37
rect 65 -41 67 -39
rect 95 -41 97 -38
rect 103 -39 113 -37
rect 103 -41 105 -39
rect 134 -41 136 -26
rect 252 -37 254 -34
rect 382 -45 384 -41
rect 390 -45 392 -41
rect 425 -43 427 -40
rect 14 -49 16 -45
rect 57 -49 59 -45
rect 65 -49 67 -45
rect 95 -49 97 -45
rect 103 -49 105 -45
rect 134 -48 136 -45
rect 198 -52 200 -49
rect 14 -74 16 -70
rect 22 -72 32 -70
rect 22 -74 24 -72
rect 57 -74 59 -70
rect 95 -74 97 -70
rect 134 -72 136 -69
rect 198 -75 200 -60
rect 382 -66 384 -53
rect 390 -63 392 -53
rect 390 -65 402 -63
rect 390 -66 392 -65
rect 400 -66 402 -65
rect 425 -66 427 -51
rect 382 -74 384 -70
rect 390 -74 392 -70
rect 425 -73 427 -70
rect 14 -87 16 -82
rect 22 -85 24 -82
rect 57 -88 59 -82
rect 95 -88 97 -82
rect 14 -95 16 -91
rect 57 -95 59 -92
rect 65 -93 75 -91
rect 65 -95 67 -93
rect 95 -95 97 -92
rect 103 -93 113 -91
rect 103 -95 105 -93
rect 134 -95 136 -80
rect 198 -82 200 -79
rect 382 -96 384 -92
rect 390 -96 392 -92
rect 425 -94 427 -91
rect 14 -103 16 -99
rect 57 -103 59 -99
rect 65 -103 67 -99
rect 95 -103 97 -99
rect 103 -103 105 -99
rect 134 -102 136 -99
rect 252 -104 254 -96
rect 252 -118 254 -112
rect 382 -117 384 -104
rect 390 -114 392 -104
rect 390 -116 402 -114
rect 390 -117 392 -116
rect 400 -117 402 -116
rect 425 -117 427 -102
rect 14 -128 16 -124
rect 22 -126 32 -124
rect 22 -128 24 -126
rect 57 -128 59 -124
rect 95 -128 97 -124
rect 134 -126 136 -123
rect 382 -125 384 -121
rect 390 -125 392 -121
rect 425 -124 427 -121
rect 14 -141 16 -136
rect 22 -139 24 -136
rect 57 -142 59 -136
rect 95 -142 97 -136
rect 14 -149 16 -145
rect 57 -149 59 -146
rect 65 -147 75 -145
rect 65 -149 67 -147
rect 95 -149 97 -146
rect 103 -147 113 -145
rect 103 -149 105 -147
rect 134 -149 136 -134
rect 252 -136 254 -130
rect 252 -148 254 -144
rect 382 -147 384 -143
rect 390 -147 392 -143
rect 425 -145 427 -142
rect 14 -157 16 -153
rect 57 -157 59 -153
rect 65 -157 67 -153
rect 95 -157 97 -153
rect 103 -157 105 -153
rect 134 -156 136 -153
rect 382 -168 384 -155
rect 390 -165 392 -155
rect 390 -167 402 -165
rect 390 -168 392 -167
rect 400 -168 402 -167
rect 425 -168 427 -153
rect 382 -176 384 -172
rect 390 -176 392 -172
rect 425 -175 427 -172
rect 14 -182 16 -178
rect 22 -180 32 -178
rect 22 -182 24 -180
rect 57 -182 59 -178
rect 95 -182 97 -178
rect 134 -180 136 -177
rect 14 -195 16 -190
rect 22 -193 24 -190
rect 57 -196 59 -190
rect 95 -196 97 -190
rect 14 -203 16 -199
rect 57 -203 59 -200
rect 65 -201 75 -199
rect 65 -203 67 -201
rect 95 -203 97 -200
rect 103 -201 113 -199
rect 103 -203 105 -201
rect 134 -203 136 -188
rect 208 -200 210 -197
rect 14 -211 16 -207
rect 57 -211 59 -207
rect 65 -211 67 -207
rect 95 -211 97 -207
rect 103 -211 105 -207
rect 134 -210 136 -207
rect 252 -204 254 -197
rect 382 -198 384 -194
rect 390 -198 392 -194
rect 425 -196 427 -193
rect 208 -223 210 -208
rect 252 -218 254 -212
rect 382 -219 384 -206
rect 390 -216 392 -206
rect 390 -218 402 -216
rect 390 -219 392 -218
rect 400 -219 402 -218
rect 425 -219 427 -204
rect 382 -227 384 -223
rect 390 -227 392 -223
rect 425 -226 427 -223
rect 208 -230 210 -227
rect 252 -236 254 -230
rect 15 -252 17 -248
rect 23 -250 33 -248
rect 23 -252 25 -250
rect 58 -252 60 -248
rect 96 -252 98 -248
rect 135 -250 137 -247
rect 252 -248 254 -244
rect 382 -249 384 -245
rect 390 -249 392 -245
rect 425 -247 427 -244
rect 15 -265 17 -260
rect 23 -263 25 -260
rect 58 -266 60 -260
rect 96 -266 98 -260
rect 15 -273 17 -269
rect 58 -273 60 -270
rect 66 -271 76 -269
rect 66 -273 68 -271
rect 96 -273 98 -270
rect 104 -271 114 -269
rect 104 -273 106 -271
rect 135 -273 137 -258
rect 382 -270 384 -257
rect 390 -267 392 -257
rect 390 -269 402 -267
rect 390 -270 392 -269
rect 400 -270 402 -269
rect 425 -270 427 -255
rect 15 -281 17 -277
rect 58 -281 60 -277
rect 66 -281 68 -277
rect 96 -281 98 -277
rect 104 -281 106 -277
rect 135 -280 137 -277
rect 382 -278 384 -274
rect 390 -278 392 -274
rect 425 -277 427 -274
rect 15 -306 17 -302
rect 23 -304 33 -302
rect 23 -306 25 -304
rect 58 -306 60 -302
rect 96 -306 98 -302
rect 135 -304 137 -301
rect 15 -319 17 -314
rect 23 -317 25 -314
rect 58 -320 60 -314
rect 96 -320 98 -314
rect 15 -327 17 -323
rect 58 -327 60 -324
rect 66 -325 76 -323
rect 66 -327 68 -325
rect 96 -327 98 -324
rect 104 -325 114 -323
rect 104 -327 106 -325
rect 135 -327 137 -312
rect 252 -314 254 -307
rect 252 -328 254 -322
rect 15 -335 17 -331
rect 58 -335 60 -331
rect 66 -335 68 -331
rect 96 -335 98 -331
rect 104 -335 106 -331
rect 135 -334 137 -331
rect 252 -346 254 -340
rect 15 -360 17 -356
rect 23 -358 33 -356
rect 23 -360 25 -358
rect 58 -360 60 -356
rect 96 -360 98 -356
rect 135 -358 137 -355
rect 252 -358 254 -354
rect 15 -373 17 -368
rect 23 -371 25 -368
rect 58 -374 60 -368
rect 96 -374 98 -368
rect 15 -381 17 -377
rect 58 -381 60 -378
rect 66 -379 76 -377
rect 66 -381 68 -379
rect 96 -381 98 -378
rect 104 -379 114 -377
rect 104 -381 106 -379
rect 135 -381 137 -366
rect 15 -389 17 -385
rect 58 -389 60 -385
rect 66 -389 68 -385
rect 96 -389 98 -385
rect 104 -389 106 -385
rect 135 -388 137 -385
rect 252 -397 254 -390
rect 15 -414 17 -410
rect 23 -412 33 -410
rect 23 -414 25 -412
rect 58 -414 60 -410
rect 96 -414 98 -410
rect 135 -412 137 -409
rect 252 -411 254 -405
rect 15 -427 17 -422
rect 23 -425 25 -422
rect 58 -428 60 -422
rect 96 -428 98 -422
rect 15 -435 17 -431
rect 58 -435 60 -432
rect 66 -433 76 -431
rect 66 -435 68 -433
rect 96 -435 98 -432
rect 104 -433 114 -431
rect 104 -435 106 -433
rect 135 -435 137 -420
rect 252 -429 254 -423
rect 15 -443 17 -439
rect 58 -443 60 -439
rect 66 -443 68 -439
rect 96 -443 98 -439
rect 104 -443 106 -439
rect 135 -442 137 -439
rect 252 -440 254 -437
rect 198 -455 200 -452
rect 15 -468 17 -464
rect 23 -466 33 -464
rect 23 -468 25 -466
rect 58 -468 60 -464
rect 96 -468 98 -464
rect 135 -466 137 -463
rect 15 -481 17 -476
rect 23 -479 25 -476
rect 58 -482 60 -476
rect 96 -482 98 -476
rect 15 -489 17 -485
rect 58 -489 60 -486
rect 66 -487 76 -485
rect 66 -489 68 -487
rect 96 -489 98 -486
rect 104 -487 114 -485
rect 104 -489 106 -487
rect 135 -489 137 -474
rect 198 -478 200 -463
rect 198 -485 200 -482
rect 15 -497 17 -493
rect 58 -497 60 -493
rect 66 -497 68 -493
rect 96 -497 98 -493
rect 104 -497 106 -493
rect 135 -496 137 -493
rect 252 -507 254 -499
rect 252 -521 254 -515
rect 252 -539 254 -533
rect 252 -551 254 -547
rect 208 -603 210 -600
rect 252 -607 254 -600
rect 208 -626 210 -611
rect 252 -621 254 -615
rect 208 -633 210 -630
rect 252 -639 254 -633
rect 252 -651 254 -647
rect 252 -717 254 -710
rect 252 -731 254 -725
rect 252 -749 254 -743
rect 252 -761 254 -757
rect 252 -802 254 -795
rect 252 -816 254 -810
rect 252 -834 254 -828
rect 252 -845 254 -842
rect 198 -860 200 -857
rect 198 -883 200 -868
rect 198 -890 200 -887
rect 252 -912 254 -904
rect 252 -926 254 -920
rect 252 -944 254 -938
rect 252 -956 254 -952
rect 208 -1008 210 -1005
rect 252 -1012 254 -1005
rect 208 -1031 210 -1016
rect 252 -1026 254 -1020
rect 208 -1038 210 -1035
rect 252 -1044 254 -1038
rect 252 -1056 254 -1052
rect 252 -1122 254 -1115
rect 252 -1136 254 -1130
rect 252 -1154 254 -1148
rect 252 -1166 254 -1162
<< polycontact >>
rect 250 833 254 837
rect 250 779 254 783
rect 193 748 197 752
rect 250 724 254 728
rect 250 668 254 672
rect 250 623 254 627
rect 203 600 207 604
rect 250 568 254 572
rect 250 513 254 517
rect 250 458 254 462
rect 250 421 254 425
rect 250 367 254 371
rect 193 336 197 340
rect 250 312 254 316
rect 250 256 254 260
rect 250 211 254 215
rect 203 188 207 192
rect 250 156 254 160
rect 250 101 254 105
rect 250 46 254 50
rect 32 34 36 38
rect 12 17 16 21
rect 55 16 59 20
rect 75 13 79 17
rect 93 16 97 20
rect 130 16 134 20
rect 251 13 255 17
rect 32 -20 36 -16
rect 12 -37 16 -33
rect 55 -38 59 -34
rect 75 -41 79 -37
rect 93 -38 97 -34
rect 130 -38 134 -34
rect 251 -41 255 -37
rect 32 -74 36 -70
rect 194 -72 198 -68
rect 378 -63 382 -59
rect 421 -63 425 -59
rect 400 -70 404 -66
rect 12 -91 16 -87
rect 55 -92 59 -88
rect 75 -95 79 -91
rect 93 -92 97 -88
rect 130 -92 134 -88
rect 251 -96 255 -92
rect 378 -114 382 -110
rect 421 -114 425 -110
rect 400 -121 404 -117
rect 32 -128 36 -124
rect 12 -145 16 -141
rect 55 -146 59 -142
rect 75 -149 79 -145
rect 93 -146 97 -142
rect 130 -146 134 -142
rect 251 -152 255 -148
rect 378 -165 382 -161
rect 421 -165 425 -161
rect 400 -172 404 -168
rect 32 -182 36 -178
rect 12 -199 16 -195
rect 55 -200 59 -196
rect 75 -203 79 -199
rect 93 -200 97 -196
rect 130 -200 134 -196
rect 251 -197 255 -193
rect 204 -220 208 -216
rect 378 -216 382 -212
rect 421 -216 425 -212
rect 400 -223 404 -219
rect 33 -252 37 -248
rect 251 -252 255 -248
rect 13 -269 17 -265
rect 56 -270 60 -266
rect 76 -273 80 -269
rect 94 -270 98 -266
rect 131 -270 135 -266
rect 378 -267 382 -263
rect 421 -267 425 -263
rect 400 -274 404 -270
rect 33 -306 37 -302
rect 251 -307 255 -303
rect 13 -323 17 -319
rect 56 -324 60 -320
rect 76 -327 80 -323
rect 94 -324 98 -320
rect 131 -324 135 -320
rect 33 -360 37 -356
rect 251 -362 255 -358
rect 13 -377 17 -373
rect 56 -378 60 -374
rect 76 -381 80 -377
rect 94 -378 98 -374
rect 131 -378 135 -374
rect 251 -390 255 -386
rect 33 -414 37 -410
rect 13 -431 17 -427
rect 56 -432 60 -428
rect 76 -435 80 -431
rect 94 -432 98 -428
rect 131 -432 135 -428
rect 251 -444 255 -440
rect 33 -468 37 -464
rect 13 -485 17 -481
rect 56 -486 60 -482
rect 76 -489 80 -485
rect 94 -486 98 -482
rect 131 -486 135 -482
rect 194 -475 198 -471
rect 251 -499 255 -495
rect 251 -555 255 -551
rect 251 -600 255 -596
rect 204 -623 208 -619
rect 251 -655 255 -651
rect 251 -710 255 -706
rect 251 -765 255 -761
rect 251 -795 255 -791
rect 251 -849 255 -845
rect 194 -880 198 -876
rect 251 -904 255 -900
rect 251 -960 255 -956
rect 251 -1005 255 -1001
rect 204 -1028 208 -1024
rect 251 -1060 255 -1056
rect 251 -1115 255 -1111
rect 251 -1170 255 -1166
<< metal1 >>
rect 250 837 254 842
rect 232 818 246 826
rect 258 818 272 826
rect 232 794 239 818
rect 258 803 262 810
rect 265 808 272 818
rect 265 794 272 801
rect 232 786 246 794
rect 258 786 272 794
rect 189 772 210 776
rect 192 768 196 772
rect 200 752 204 760
rect 232 754 239 786
rect 215 752 239 754
rect 186 748 193 752
rect 200 748 239 752
rect 200 745 204 748
rect 215 747 239 748
rect 192 737 196 741
rect 185 733 202 737
rect 209 733 210 737
rect 232 716 239 747
rect 250 744 254 779
rect 250 728 254 739
rect 232 708 246 716
rect 258 708 305 716
rect 232 684 239 708
rect 258 693 262 700
rect 265 684 272 708
rect 232 676 246 684
rect 258 676 272 684
rect 250 656 254 668
rect 150 650 249 654
rect 150 456 154 650
rect 186 604 192 650
rect 195 624 215 628
rect 250 627 254 649
rect 202 620 206 624
rect 265 622 272 676
rect 264 616 272 622
rect 210 604 214 612
rect 232 608 246 616
rect 258 608 272 616
rect 186 600 203 604
rect 210 600 219 604
rect 210 597 214 600
rect 202 589 206 593
rect 194 588 220 589
rect 201 585 220 588
rect 232 584 239 608
rect 257 593 261 600
rect 264 597 272 608
rect 265 584 272 597
rect 232 576 246 584
rect 258 576 272 584
rect 232 543 239 576
rect 217 537 232 543
rect 211 536 232 537
rect 232 506 239 536
rect 250 564 254 568
rect 250 517 254 559
rect 232 498 246 506
rect 258 498 272 506
rect 232 474 239 498
rect 258 483 262 490
rect 265 488 272 498
rect 265 474 272 481
rect 232 466 246 474
rect 258 466 272 474
rect 250 456 254 458
rect 149 452 254 456
rect 4 44 94 45
rect 4 41 147 44
rect 9 34 13 41
rect 5 17 12 21
rect 25 13 29 26
rect 37 20 41 33
rect 52 34 56 41
rect 90 40 147 41
rect 90 34 94 40
rect 129 36 133 40
rect 64 26 82 30
rect 102 26 124 30
rect 37 16 55 20
rect 68 13 72 26
rect 78 23 82 26
rect 78 20 88 23
rect 21 9 37 13
rect 9 4 13 9
rect 84 16 93 20
rect 106 13 110 26
rect 121 20 124 26
rect 137 20 141 28
rect 150 20 154 452
rect 250 425 254 429
rect 232 406 246 414
rect 258 406 272 414
rect 232 382 239 406
rect 258 391 262 398
rect 265 396 272 406
rect 265 382 272 389
rect 232 374 246 382
rect 258 374 272 382
rect 189 360 210 364
rect 192 356 196 360
rect 200 340 204 348
rect 232 342 239 374
rect 215 340 239 342
rect 185 336 193 340
rect 200 336 239 340
rect 200 333 204 336
rect 215 335 239 336
rect 192 325 196 329
rect 185 321 201 325
rect 208 321 210 325
rect 232 304 239 335
rect 250 332 254 367
rect 250 316 254 327
rect 232 296 246 304
rect 258 296 305 304
rect 232 272 239 296
rect 258 281 262 288
rect 265 272 272 296
rect 232 264 246 272
rect 258 264 272 272
rect 250 244 254 256
rect 121 16 130 20
rect 137 16 154 20
rect 157 238 249 242
rect 157 44 161 238
rect 188 192 192 238
rect 195 212 212 216
rect 217 212 220 216
rect 250 215 254 237
rect 202 208 206 212
rect 265 210 272 264
rect 264 204 272 210
rect 210 192 214 200
rect 232 196 246 204
rect 258 196 272 204
rect 188 188 203 192
rect 210 188 219 192
rect 210 185 214 188
rect 202 177 206 181
rect 195 176 220 177
rect 195 173 203 176
rect 208 173 220 176
rect 232 172 239 196
rect 257 181 261 188
rect 264 185 272 196
rect 265 172 272 185
rect 232 164 246 172
rect 258 164 272 172
rect 232 131 239 164
rect 215 129 232 131
rect 219 124 232 129
rect 232 94 239 124
rect 250 152 254 156
rect 250 105 254 147
rect 232 86 246 94
rect 258 86 272 94
rect 232 62 239 86
rect 258 71 262 78
rect 265 76 272 86
rect 265 62 272 69
rect 232 54 246 62
rect 258 54 272 62
rect 250 44 254 46
rect 157 40 254 44
rect 137 13 141 16
rect 52 4 56 9
rect 90 5 94 9
rect 129 5 133 9
rect 90 4 147 5
rect -9 0 147 4
rect -9 -50 -5 0
rect 4 -10 94 -9
rect 4 -13 147 -10
rect 9 -20 13 -13
rect 5 -37 12 -33
rect 25 -41 29 -28
rect 37 -34 41 -21
rect 52 -20 56 -13
rect 90 -14 147 -13
rect 90 -20 94 -14
rect 129 -18 133 -14
rect 64 -28 82 -24
rect 102 -28 124 -24
rect 37 -38 55 -34
rect 68 -41 72 -28
rect 78 -31 82 -28
rect 78 -34 88 -31
rect 21 -45 37 -41
rect 9 -50 13 -45
rect 84 -38 93 -34
rect 106 -41 110 -28
rect 121 -34 124 -28
rect 137 -34 141 -26
rect 157 -34 161 40
rect 251 17 255 22
rect 121 -38 130 -34
rect 137 -38 161 -34
rect 233 -2 247 6
rect 259 -2 273 6
rect 233 -26 240 -2
rect 259 -17 263 -10
rect 266 -12 273 -2
rect 266 -26 273 -19
rect 233 -34 247 -26
rect 259 -34 273 -26
rect 137 -41 141 -38
rect 52 -50 56 -45
rect 90 -49 94 -45
rect 129 -49 133 -45
rect 186 -48 206 -43
rect 90 -50 147 -49
rect -9 -54 147 -50
rect 193 -52 197 -48
rect -9 -104 -5 -54
rect 4 -64 94 -63
rect 4 -67 147 -64
rect 9 -74 13 -67
rect 5 -91 12 -87
rect 25 -95 29 -82
rect 37 -88 41 -75
rect 52 -74 56 -67
rect 90 -68 147 -67
rect 201 -68 205 -60
rect 233 -66 240 -34
rect 216 -68 240 -66
rect 90 -74 94 -68
rect 129 -72 133 -68
rect 64 -82 82 -78
rect 102 -82 124 -78
rect 187 -72 194 -68
rect 201 -72 240 -68
rect 201 -75 205 -72
rect 216 -73 240 -72
rect 37 -92 55 -88
rect 68 -95 72 -82
rect 78 -85 82 -82
rect 78 -88 88 -85
rect 21 -99 37 -95
rect 9 -104 13 -99
rect 84 -92 93 -88
rect 106 -95 110 -82
rect 121 -88 124 -82
rect 137 -88 141 -80
rect 193 -83 197 -79
rect 186 -87 202 -83
rect 121 -92 130 -88
rect 137 -92 175 -88
rect 209 -87 211 -83
rect 137 -95 141 -92
rect 52 -104 56 -99
rect 90 -103 94 -99
rect 129 -103 133 -99
rect 90 -104 147 -103
rect -9 -108 147 -104
rect -9 -158 -5 -108
rect 4 -118 94 -117
rect 4 -121 147 -118
rect 9 -128 13 -121
rect 5 -145 12 -141
rect 25 -149 29 -136
rect 37 -142 41 -129
rect 52 -128 56 -121
rect 90 -122 147 -121
rect 90 -128 94 -122
rect 129 -126 133 -122
rect 64 -136 82 -132
rect 102 -136 124 -132
rect 37 -146 55 -142
rect 68 -149 72 -136
rect 78 -139 82 -136
rect 78 -142 88 -139
rect 21 -153 37 -149
rect 9 -158 13 -153
rect 84 -146 93 -142
rect 106 -149 110 -136
rect 121 -142 124 -136
rect 137 -142 141 -134
rect 121 -146 130 -142
rect 137 -146 160 -142
rect 137 -149 141 -146
rect 52 -158 56 -153
rect 90 -157 94 -153
rect 129 -157 133 -153
rect 90 -158 147 -157
rect -9 -162 147 -158
rect -9 -212 -5 -162
rect 4 -172 94 -171
rect 4 -175 147 -172
rect 9 -182 13 -175
rect 5 -199 12 -195
rect 25 -203 29 -190
rect 37 -196 41 -183
rect 52 -182 56 -175
rect 90 -176 147 -175
rect 90 -182 94 -176
rect 129 -180 133 -176
rect 64 -190 82 -186
rect 102 -190 124 -186
rect 37 -200 55 -196
rect 68 -203 72 -190
rect 78 -193 82 -190
rect 78 -196 88 -193
rect 21 -207 37 -203
rect 9 -212 13 -207
rect 84 -200 93 -196
rect 106 -203 110 -190
rect 121 -196 124 -190
rect 137 -196 141 -188
rect 121 -200 130 -196
rect 137 -200 153 -196
rect 137 -203 141 -200
rect 52 -212 56 -207
rect 90 -211 94 -207
rect 129 -211 133 -207
rect 90 -212 147 -211
rect -9 -216 147 -212
rect -9 -282 -5 -216
rect 150 -223 153 -200
rect 146 -226 153 -223
rect 5 -242 95 -241
rect 5 -245 148 -242
rect 10 -252 14 -245
rect 6 -269 13 -265
rect 26 -273 30 -260
rect 38 -266 42 -253
rect 53 -252 57 -245
rect 91 -246 148 -245
rect 91 -252 95 -246
rect 130 -250 134 -246
rect 65 -260 83 -256
rect 103 -260 125 -256
rect 38 -270 56 -266
rect 69 -273 73 -260
rect 79 -263 83 -260
rect 79 -266 89 -263
rect 22 -277 38 -273
rect 10 -282 14 -277
rect 85 -270 94 -266
rect 107 -273 111 -260
rect 122 -266 125 -260
rect 138 -266 142 -258
rect 156 -257 160 -146
rect 171 -166 175 -92
rect 233 -104 240 -73
rect 376 -38 438 -34
rect 251 -76 255 -41
rect 377 -45 381 -38
rect 393 -45 397 -38
rect 420 -43 424 -38
rect 385 -59 389 -53
rect 428 -59 432 -51
rect 377 -63 378 -59
rect 385 -63 421 -59
rect 428 -63 441 -59
rect 393 -66 397 -63
rect 428 -66 432 -63
rect 404 -70 405 -66
rect 377 -75 381 -70
rect 420 -74 424 -70
rect 413 -75 438 -74
rect 364 -79 438 -75
rect 251 -92 255 -81
rect 233 -112 247 -104
rect 259 -112 306 -104
rect 233 -136 240 -112
rect 259 -127 263 -120
rect 266 -136 273 -112
rect 233 -144 247 -136
rect 259 -144 273 -136
rect 251 -164 255 -152
rect 171 -170 250 -166
rect 156 -261 164 -257
rect 122 -270 131 -266
rect 138 -270 151 -266
rect 138 -273 142 -270
rect 53 -282 57 -277
rect 91 -281 95 -277
rect 130 -281 134 -277
rect 91 -282 148 -281
rect -9 -286 148 -282
rect -9 -336 -5 -286
rect 5 -296 95 -295
rect 5 -299 148 -296
rect 10 -306 14 -299
rect 6 -323 13 -319
rect 26 -327 30 -314
rect 38 -320 42 -307
rect 53 -306 57 -299
rect 91 -300 148 -299
rect 91 -306 95 -300
rect 130 -304 134 -300
rect 65 -314 83 -310
rect 103 -314 125 -310
rect 38 -324 56 -320
rect 69 -327 73 -314
rect 79 -317 83 -314
rect 79 -320 89 -317
rect 22 -331 38 -327
rect 10 -336 14 -331
rect 85 -324 94 -320
rect 107 -327 111 -314
rect 122 -320 125 -314
rect 138 -320 142 -312
rect 122 -324 131 -320
rect 138 -324 151 -320
rect 138 -327 142 -324
rect 53 -336 57 -331
rect 91 -335 95 -331
rect 130 -335 134 -331
rect 91 -336 148 -335
rect -9 -340 148 -336
rect -9 -390 -5 -340
rect 5 -350 95 -349
rect 5 -353 148 -350
rect 10 -360 14 -353
rect 6 -377 13 -373
rect 26 -381 30 -368
rect 38 -374 42 -361
rect 53 -360 57 -353
rect 91 -354 148 -353
rect 91 -360 95 -354
rect 130 -358 134 -354
rect 65 -368 83 -364
rect 103 -368 125 -364
rect 38 -378 56 -374
rect 69 -381 73 -368
rect 79 -371 83 -368
rect 79 -374 89 -371
rect 22 -385 38 -381
rect 10 -390 14 -385
rect 85 -378 94 -374
rect 107 -381 111 -368
rect 122 -374 125 -368
rect 138 -374 142 -366
rect 122 -378 131 -374
rect 138 -378 151 -374
rect 138 -381 142 -378
rect 53 -390 57 -385
rect 91 -389 95 -385
rect 130 -389 134 -385
rect 91 -390 148 -389
rect -9 -394 148 -390
rect -9 -444 -5 -394
rect 5 -404 95 -403
rect 5 -407 148 -404
rect 10 -414 14 -407
rect 6 -431 13 -427
rect 26 -435 30 -422
rect 38 -428 42 -415
rect 53 -414 57 -407
rect 91 -408 148 -407
rect 91 -414 95 -408
rect 130 -412 134 -408
rect 65 -422 83 -418
rect 103 -422 125 -418
rect 38 -432 56 -428
rect 69 -435 73 -422
rect 79 -425 83 -422
rect 79 -428 89 -425
rect 22 -439 38 -435
rect 10 -444 14 -439
rect 85 -432 94 -428
rect 107 -435 111 -422
rect 122 -428 125 -422
rect 138 -428 142 -420
rect 122 -432 131 -428
rect 138 -432 151 -428
rect 138 -435 142 -432
rect 53 -444 57 -439
rect 91 -443 95 -439
rect 130 -443 134 -439
rect 91 -444 148 -443
rect -9 -448 148 -444
rect -9 -498 -5 -448
rect 5 -458 95 -457
rect 5 -461 148 -458
rect 10 -468 14 -461
rect 6 -485 13 -481
rect 26 -489 30 -476
rect 38 -482 42 -469
rect 53 -468 57 -461
rect 91 -462 148 -461
rect 91 -468 95 -462
rect 130 -466 134 -462
rect 65 -476 83 -472
rect 103 -476 125 -472
rect 38 -486 56 -482
rect 69 -489 73 -476
rect 79 -479 83 -476
rect 79 -482 89 -479
rect 22 -493 38 -489
rect 10 -498 14 -493
rect 85 -486 94 -482
rect 107 -489 111 -476
rect 122 -482 125 -476
rect 138 -482 142 -474
rect 122 -486 131 -482
rect 138 -486 155 -482
rect 138 -489 142 -486
rect 53 -498 57 -493
rect 91 -497 95 -493
rect 130 -497 134 -493
rect 91 -498 148 -497
rect -9 -502 148 -498
rect 131 -1183 135 -502
rect 151 -876 155 -486
rect 160 -569 164 -261
rect 178 -366 182 -170
rect 189 -216 193 -170
rect 196 -196 213 -192
rect 218 -196 221 -192
rect 251 -193 255 -172
rect 203 -200 207 -196
rect 266 -198 273 -144
rect 265 -204 273 -198
rect 211 -216 215 -208
rect 233 -212 247 -204
rect 259 -212 273 -204
rect 189 -220 204 -216
rect 211 -220 220 -216
rect 211 -223 215 -220
rect 203 -231 207 -227
rect 196 -235 213 -231
rect 233 -236 240 -212
rect 258 -227 262 -220
rect 265 -223 273 -212
rect 266 -236 273 -223
rect 233 -244 247 -236
rect 259 -244 273 -236
rect 364 -126 368 -79
rect 377 -89 438 -85
rect 377 -96 381 -89
rect 393 -96 397 -89
rect 420 -94 424 -89
rect 385 -110 389 -104
rect 428 -110 432 -102
rect 377 -114 378 -110
rect 385 -114 421 -110
rect 428 -114 441 -110
rect 393 -117 397 -114
rect 428 -117 432 -114
rect 377 -126 381 -121
rect 420 -125 424 -121
rect 413 -126 438 -125
rect 364 -130 438 -126
rect 364 -177 368 -130
rect 377 -140 438 -136
rect 377 -147 381 -140
rect 393 -147 397 -140
rect 420 -145 424 -140
rect 385 -161 389 -155
rect 428 -161 432 -153
rect 385 -165 421 -161
rect 428 -165 441 -161
rect 393 -168 397 -165
rect 428 -168 432 -165
rect 404 -169 409 -168
rect 377 -177 381 -172
rect 420 -176 424 -172
rect 413 -177 438 -176
rect 364 -181 438 -177
rect 364 -228 368 -181
rect 377 -191 438 -187
rect 377 -198 381 -191
rect 393 -198 397 -191
rect 420 -196 424 -191
rect 385 -212 389 -206
rect 428 -212 432 -204
rect 385 -216 421 -212
rect 428 -216 441 -212
rect 393 -219 397 -216
rect 428 -219 432 -216
rect 377 -228 381 -223
rect 420 -227 424 -223
rect 413 -228 438 -227
rect 364 -232 438 -228
rect 233 -277 240 -244
rect 220 -284 233 -277
rect 233 -314 240 -284
rect 251 -256 255 -252
rect 251 -303 255 -261
rect 364 -279 368 -232
rect 377 -242 438 -238
rect 377 -249 381 -242
rect 393 -249 397 -242
rect 420 -247 424 -242
rect 385 -263 389 -257
rect 428 -263 432 -255
rect 385 -267 421 -263
rect 428 -267 441 -263
rect 393 -270 397 -267
rect 428 -270 432 -267
rect 377 -279 381 -274
rect 420 -278 424 -274
rect 413 -279 438 -278
rect 364 -283 438 -279
rect 233 -322 247 -314
rect 259 -322 273 -314
rect 233 -346 240 -322
rect 259 -337 263 -330
rect 266 -332 273 -322
rect 266 -346 273 -339
rect 233 -354 247 -346
rect 259 -354 273 -346
rect 251 -366 255 -362
rect 178 -370 255 -366
rect 251 -386 255 -381
rect 233 -405 247 -397
rect 259 -405 273 -397
rect 233 -429 240 -405
rect 259 -420 263 -413
rect 266 -415 273 -405
rect 266 -429 273 -422
rect 233 -437 247 -429
rect 259 -437 273 -429
rect 186 -450 189 -447
rect 194 -450 211 -447
rect 186 -451 211 -450
rect 193 -455 197 -451
rect 201 -471 205 -463
rect 233 -469 240 -437
rect 216 -471 240 -469
rect 187 -475 194 -471
rect 201 -475 240 -471
rect 201 -478 205 -475
rect 216 -476 240 -475
rect 193 -486 197 -482
rect 186 -490 201 -486
rect 209 -490 211 -486
rect 233 -507 240 -476
rect 251 -479 255 -444
rect 251 -495 255 -484
rect 233 -515 247 -507
rect 259 -515 306 -507
rect 233 -539 240 -515
rect 259 -530 263 -523
rect 266 -539 273 -515
rect 233 -547 247 -539
rect 259 -547 273 -539
rect 251 -568 255 -555
rect 160 -573 251 -569
rect 160 -619 164 -573
rect 196 -599 213 -595
rect 203 -603 207 -599
rect 218 -599 221 -595
rect 251 -596 255 -573
rect 266 -601 273 -547
rect 265 -607 273 -601
rect 211 -619 215 -611
rect 233 -615 247 -607
rect 259 -615 273 -607
rect 160 -623 204 -619
rect 211 -623 220 -619
rect 185 -769 189 -623
rect 211 -626 215 -623
rect 203 -634 207 -630
rect 196 -638 214 -634
rect 233 -639 240 -615
rect 258 -630 262 -623
rect 265 -626 273 -615
rect 266 -639 273 -626
rect 233 -647 247 -639
rect 259 -647 273 -639
rect 233 -680 240 -647
rect 221 -687 233 -680
rect 233 -717 240 -687
rect 251 -659 255 -655
rect 251 -706 255 -664
rect 233 -725 247 -717
rect 259 -725 273 -717
rect 233 -749 240 -725
rect 259 -740 263 -733
rect 266 -735 273 -725
rect 266 -749 273 -742
rect 233 -757 247 -749
rect 259 -757 273 -749
rect 251 -769 255 -765
rect 185 -773 255 -769
rect 254 -785 255 -783
rect 251 -791 255 -785
rect 233 -810 247 -802
rect 259 -810 273 -802
rect 233 -834 240 -810
rect 259 -825 263 -818
rect 266 -820 273 -810
rect 266 -834 273 -827
rect 233 -842 247 -834
rect 259 -842 273 -834
rect 186 -855 190 -852
rect 195 -855 211 -852
rect 186 -856 211 -855
rect 193 -860 197 -856
rect 201 -876 205 -868
rect 233 -874 240 -842
rect 216 -876 240 -874
rect 151 -880 194 -876
rect 201 -880 240 -876
rect 151 -974 155 -880
rect 201 -883 205 -880
rect 216 -881 240 -880
rect 193 -891 197 -887
rect 189 -895 211 -891
rect 233 -912 240 -881
rect 251 -884 255 -849
rect 251 -900 255 -889
rect 233 -920 247 -912
rect 259 -920 306 -912
rect 233 -944 240 -920
rect 259 -935 263 -928
rect 266 -944 273 -920
rect 233 -952 247 -944
rect 259 -952 273 -944
rect 251 -972 255 -960
rect 151 -978 250 -974
rect 152 -1172 156 -978
rect 196 -1003 214 -1000
rect 219 -1003 221 -1000
rect 196 -1004 221 -1003
rect 251 -1001 255 -979
rect 203 -1008 207 -1004
rect 266 -1006 273 -952
rect 265 -1012 273 -1006
rect 211 -1024 215 -1016
rect 233 -1020 247 -1012
rect 259 -1020 273 -1012
rect 198 -1028 204 -1024
rect 211 -1028 220 -1024
rect 211 -1031 215 -1028
rect 203 -1039 207 -1035
rect 196 -1043 221 -1039
rect 196 -1053 200 -1043
rect 233 -1044 240 -1020
rect 258 -1035 262 -1028
rect 265 -1031 273 -1020
rect 266 -1044 273 -1031
rect 233 -1052 247 -1044
rect 259 -1052 273 -1044
rect 233 -1085 240 -1052
rect 216 -1088 233 -1085
rect 216 -1089 217 -1088
rect 214 -1092 217 -1089
rect 224 -1092 233 -1088
rect 233 -1122 240 -1092
rect 251 -1064 255 -1060
rect 251 -1111 255 -1069
rect 233 -1130 247 -1122
rect 259 -1130 273 -1122
rect 233 -1154 240 -1130
rect 259 -1145 263 -1138
rect 266 -1140 273 -1130
rect 266 -1154 273 -1147
rect 233 -1162 247 -1154
rect 259 -1162 273 -1154
rect 251 -1172 255 -1170
rect 152 -1176 255 -1172
rect 364 -1183 368 -283
rect 131 -1187 368 -1183
<< m2contact >>
rect 265 801 272 808
rect 184 772 189 777
rect 181 748 186 753
rect 250 739 255 744
rect 215 624 220 629
rect 219 600 224 605
rect 211 537 217 543
rect 250 559 255 564
rect 265 481 272 488
rect -1 41 4 46
rect 36 33 41 38
rect 37 8 42 13
rect 250 429 255 434
rect 265 389 272 396
rect 184 360 189 365
rect 179 334 185 340
rect 250 327 255 332
rect 212 212 217 217
rect 219 188 224 193
rect 213 124 219 129
rect 250 147 255 152
rect 265 69 272 76
rect 75 8 80 13
rect -1 -13 4 -8
rect 36 -21 41 -16
rect 37 -46 42 -41
rect 251 22 256 27
rect 266 -19 273 -12
rect 75 -46 80 -41
rect 206 -48 211 -43
rect -1 -67 4 -62
rect 36 -75 41 -70
rect 181 -73 187 -68
rect 37 -100 42 -95
rect 75 -100 80 -95
rect -1 -121 4 -116
rect 36 -129 41 -124
rect 37 -154 42 -149
rect 75 -154 80 -149
rect -1 -175 4 -170
rect 36 -183 41 -178
rect 37 -208 42 -203
rect 75 -208 80 -203
rect 0 -245 5 -240
rect 37 -253 42 -248
rect 38 -278 43 -273
rect 371 -38 376 -33
rect 251 -81 256 -76
rect 151 -270 156 -265
rect 76 -278 81 -273
rect 0 -299 5 -294
rect 37 -307 42 -302
rect 38 -332 43 -327
rect 151 -324 156 -319
rect 76 -332 81 -327
rect 0 -353 5 -348
rect 37 -361 42 -356
rect 38 -386 43 -381
rect 151 -378 156 -373
rect 76 -386 81 -381
rect 0 -407 5 -402
rect 37 -415 42 -410
rect 38 -440 43 -435
rect 151 -432 156 -427
rect 76 -440 81 -435
rect 0 -461 5 -456
rect 37 -469 42 -464
rect 38 -494 43 -489
rect 76 -494 81 -489
rect 213 -196 218 -191
rect 220 -220 225 -215
rect 372 -89 377 -84
rect 372 -140 377 -135
rect 372 -191 377 -186
rect 214 -284 220 -277
rect 251 -261 256 -256
rect 372 -242 377 -237
rect 266 -339 273 -332
rect 251 -381 256 -376
rect 266 -422 273 -415
rect 189 -450 194 -445
rect 182 -475 187 -470
rect 251 -484 256 -479
rect 213 -600 218 -595
rect 220 -623 225 -618
rect 214 -687 221 -680
rect 251 -664 256 -659
rect 266 -742 273 -735
rect 249 -785 254 -780
rect 266 -827 273 -820
rect 190 -855 195 -850
rect 251 -889 256 -884
rect 214 -1003 219 -998
rect 220 -1028 225 -1023
rect 251 -1069 256 -1064
rect 266 -1147 273 -1140
<< pm12contact >>
rect 113 15 118 20
rect 113 -39 118 -34
rect 113 -93 118 -88
rect 113 -147 118 -142
rect 113 -201 118 -196
rect 114 -271 119 -266
rect 114 -325 119 -320
rect 114 -379 119 -374
rect 114 -433 119 -428
rect 114 -487 119 -482
<< metal2 >>
rect 18 856 368 861
rect 18 52 23 856
rect 184 777 189 856
rect 151 748 181 752
rect 151 543 156 748
rect 215 670 220 856
rect 272 801 289 808
rect 179 665 220 670
rect 179 543 184 665
rect 215 629 220 665
rect 224 739 250 743
rect 224 563 228 739
rect 282 594 289 801
rect 282 587 305 594
rect 224 559 250 563
rect 151 537 211 543
rect 217 537 218 543
rect -1 47 23 52
rect 37 48 117 52
rect -1 46 4 47
rect 0 -8 4 41
rect 37 38 41 48
rect 113 20 117 48
rect 42 8 75 13
rect 0 -62 4 -13
rect 37 -6 117 -2
rect 37 -16 41 -6
rect 113 -34 117 -6
rect 42 -46 75 -41
rect 0 -116 4 -67
rect 37 -60 117 -56
rect 37 -70 41 -60
rect 113 -88 117 -60
rect 42 -100 75 -95
rect 0 -170 4 -121
rect 37 -114 117 -110
rect 37 -124 41 -114
rect 113 -142 117 -114
rect 42 -154 75 -149
rect 0 -240 4 -175
rect 37 -168 117 -164
rect 37 -178 41 -168
rect 113 -196 117 -168
rect 42 -208 75 -203
rect 38 -238 118 -234
rect 0 -294 4 -245
rect 38 -248 42 -238
rect 114 -266 118 -238
rect 151 -265 156 537
rect 179 380 184 537
rect 282 488 289 587
rect 272 481 289 488
rect 272 389 289 396
rect 179 374 217 380
rect 179 360 184 374
rect 160 336 179 340
rect 160 129 165 336
rect 212 231 217 374
rect 182 226 217 231
rect 182 141 187 226
rect 212 217 217 226
rect 224 327 250 331
rect 224 151 228 327
rect 282 182 289 389
rect 282 175 305 182
rect 224 147 250 151
rect 182 136 228 141
rect 160 124 213 129
rect 43 -278 76 -273
rect 38 -292 118 -288
rect 0 -348 4 -299
rect 38 -302 42 -292
rect 114 -320 118 -292
rect 160 -319 165 124
rect 223 -29 228 136
rect 282 76 289 175
rect 272 69 289 76
rect 273 -19 290 -12
rect 206 -34 228 -29
rect 206 -43 211 -34
rect 217 -53 223 -34
rect 213 -56 223 -53
rect 156 -324 165 -319
rect 169 -72 181 -68
rect 169 -277 174 -72
rect 213 -180 218 -56
rect 189 -185 218 -180
rect 189 -268 194 -185
rect 213 -191 218 -185
rect 225 -81 251 -77
rect 225 -257 229 -81
rect 283 -226 290 -19
rect 363 -33 368 856
rect 363 -38 371 -33
rect 363 -84 368 -38
rect 363 -89 372 -84
rect 363 -135 368 -89
rect 363 -140 372 -135
rect 363 -186 368 -140
rect 363 -191 372 -186
rect 283 -233 306 -226
rect 225 -261 251 -257
rect 189 -272 264 -268
rect 169 -284 214 -277
rect 43 -332 76 -327
rect 38 -346 118 -342
rect 0 -402 4 -353
rect 38 -356 42 -346
rect 114 -374 118 -346
rect 169 -373 174 -284
rect 259 -289 264 -272
rect 156 -378 174 -373
rect 189 -293 264 -289
rect 43 -386 76 -381
rect 38 -400 118 -396
rect 0 -456 4 -407
rect 38 -410 42 -400
rect 114 -428 118 -400
rect 156 -432 178 -427
rect 43 -440 76 -435
rect 38 -454 118 -450
rect 38 -464 42 -454
rect 114 -482 118 -454
rect 173 -471 178 -432
rect 189 -434 194 -293
rect 283 -332 290 -233
rect 363 -237 368 -191
rect 363 -242 372 -237
rect 273 -339 290 -332
rect 273 -422 290 -415
rect 189 -439 218 -434
rect 189 -445 194 -439
rect 173 -475 182 -471
rect 43 -494 76 -489
rect 173 -680 178 -475
rect 213 -585 218 -439
rect 190 -590 218 -585
rect 190 -669 195 -590
rect 213 -595 218 -590
rect 225 -484 251 -480
rect 225 -660 229 -484
rect 283 -629 290 -422
rect 283 -636 306 -629
rect 225 -664 251 -660
rect 190 -676 265 -669
rect 173 -687 214 -680
rect 259 -692 265 -676
rect 190 -699 265 -692
rect 190 -837 195 -699
rect 283 -735 290 -636
rect 273 -742 290 -735
rect 273 -827 290 -820
rect 190 -842 219 -837
rect 190 -850 195 -842
rect 214 -998 219 -842
rect 225 -889 251 -885
rect 225 -1065 229 -889
rect 283 -1034 290 -827
rect 283 -1041 306 -1034
rect 225 -1069 251 -1065
rect 283 -1140 290 -1041
rect 273 -1147 290 -1140
<< m123contact >>
rect 202 731 209 738
rect 248 842 254 847
rect 194 581 201 588
rect 249 649 256 656
rect 139 -227 146 -220
rect 232 536 239 543
rect 250 429 255 434
rect 201 318 208 325
rect 203 171 208 176
rect 249 237 256 244
rect 232 124 239 131
rect 251 22 256 27
rect 202 -90 209 -83
rect 213 -238 221 -230
rect 250 -172 257 -164
rect 372 -63 377 -58
rect 405 -72 410 -66
rect 372 -114 377 -109
rect 404 -122 409 -117
rect 373 -165 378 -160
rect 404 -174 409 -169
rect 233 -284 240 -277
rect 373 -216 378 -211
rect 404 -224 409 -219
rect 373 -267 378 -262
rect 404 -275 409 -270
rect 251 -381 256 -376
rect 201 -494 209 -486
rect 214 -640 221 -633
rect 251 -573 256 -568
rect 233 -687 240 -680
rect 249 -785 254 -780
rect 182 -896 189 -889
rect 192 -1030 198 -1024
rect 195 -1061 202 -1053
rect 250 -979 257 -972
rect 217 -1095 224 -1088
rect 233 -1092 240 -1085
<< metal3 >>
rect 248 847 255 848
rect 254 846 255 847
rect 254 842 326 846
rect 248 841 255 842
rect 322 654 326 842
rect 354 654 359 655
rect 256 650 359 654
rect 239 536 348 543
rect 249 434 256 435
rect 249 429 250 434
rect 255 433 256 434
rect 255 429 314 433
rect 249 428 256 429
rect 310 242 314 429
rect 256 238 337 242
rect 202 176 209 177
rect 202 171 203 176
rect 208 171 209 176
rect 202 170 209 171
rect 231 131 240 132
rect 231 124 232 131
rect 239 124 329 131
rect 231 123 240 124
rect 250 27 257 28
rect 250 22 251 27
rect 256 26 257 27
rect 256 22 315 26
rect 250 21 257 22
rect 311 -165 315 22
rect 323 -118 328 124
rect 333 -110 337 238
rect 341 -67 348 536
rect 354 -59 359 650
rect 354 -63 372 -59
rect 341 -72 405 -67
rect 333 -114 372 -110
rect 323 -122 404 -118
rect 335 -165 373 -161
rect 257 -169 339 -165
rect 403 -169 410 -168
rect 360 -174 404 -169
rect 409 -174 410 -169
rect 277 -179 365 -174
rect 403 -175 410 -174
rect 277 -181 331 -179
rect 146 -224 169 -221
rect 166 -1024 169 -224
rect 277 -276 284 -181
rect 232 -277 284 -276
rect 232 -284 233 -277
rect 240 -283 284 -277
rect 310 -216 373 -212
rect 378 -216 382 -212
rect 240 -284 241 -283
rect 232 -285 241 -284
rect 250 -376 257 -375
rect 310 -376 315 -216
rect 250 -381 251 -376
rect 256 -381 315 -376
rect 250 -382 257 -381
rect 250 -568 257 -567
rect 310 -568 315 -381
rect 250 -573 251 -568
rect 256 -573 315 -568
rect 319 -224 404 -221
rect 250 -574 257 -573
rect 319 -679 322 -224
rect 232 -680 322 -679
rect 232 -687 233 -680
rect 240 -686 322 -680
rect 240 -687 241 -686
rect 319 -687 322 -686
rect 335 -267 373 -263
rect 232 -688 241 -687
rect 248 -780 255 -779
rect 248 -785 249 -780
rect 254 -781 255 -780
rect 254 -785 320 -781
rect 248 -786 255 -785
rect 316 -973 320 -785
rect 335 -973 339 -267
rect 257 -977 339 -973
rect 351 -275 404 -271
rect 166 -1028 192 -1024
rect 166 -1090 169 -1028
rect 166 -1093 217 -1090
rect 351 -1086 357 -275
rect 240 -1092 357 -1086
<< labels >>
rlabel metal1 -1 41 35 45 5 vdd
rlabel metal1 5 17 16 21 1 D
rlabel metal1 -1 41 94 45 1 vdd
rlabel metal1 146 3 146 3 8 gnd
rlabel metal1 90 40 147 44 1 vdd
rlabel metal1 90 0 147 5 1 gnd
rlabel metal1 -1 -54 35 -50 1 gnd
rlabel metal1 -1 -13 35 -9 5 vdd
rlabel metal1 5 -37 16 -33 1 D
rlabel metal1 -1 -54 94 -50 1 gnd
rlabel metal1 -1 -13 94 -9 1 vdd
rlabel metal1 146 -51 146 -51 8 gnd
rlabel metal1 90 -14 147 -10 1 vdd
rlabel metal1 90 -54 147 -49 1 gnd
rlabel metal1 -1 -108 35 -104 1 gnd
rlabel metal1 -1 -67 35 -63 5 vdd
rlabel metal1 5 -91 16 -87 1 D
rlabel metal1 -1 -108 94 -104 1 gnd
rlabel metal1 -1 -67 94 -63 1 vdd
rlabel metal1 146 -105 146 -105 8 gnd
rlabel metal1 90 -68 147 -64 1 vdd
rlabel metal1 90 -108 147 -103 1 gnd
rlabel metal1 -1 -162 35 -158 1 gnd
rlabel metal1 -1 -121 35 -117 5 vdd
rlabel metal1 5 -145 16 -141 1 D
rlabel metal1 -1 -162 94 -158 1 gnd
rlabel metal1 -1 -121 94 -117 1 vdd
rlabel metal1 146 -159 146 -159 8 gnd
rlabel metal1 90 -122 147 -118 1 vdd
rlabel metal1 90 -162 147 -157 1 gnd
rlabel metal1 -1 -216 35 -212 1 gnd
rlabel metal1 -1 -175 35 -171 5 vdd
rlabel metal1 5 -199 16 -195 1 D
rlabel metal1 -1 -216 94 -212 1 gnd
rlabel metal1 -1 -175 94 -171 1 vdd
rlabel metal1 90 -176 147 -172 1 vdd
rlabel metal1 0 -286 36 -282 1 gnd
rlabel metal1 0 -245 36 -241 5 vdd
rlabel metal1 6 -269 17 -265 1 D
rlabel metal1 0 -286 95 -282 1 gnd
rlabel metal1 0 -245 95 -241 1 vdd
rlabel metal1 147 -283 147 -283 8 gnd
rlabel metal1 91 -246 148 -242 1 vdd
rlabel metal1 91 -286 148 -281 1 gnd
rlabel metal1 0 -340 36 -336 1 gnd
rlabel metal1 0 -299 36 -295 5 vdd
rlabel metal1 6 -323 17 -319 1 D
rlabel metal1 0 -340 95 -336 1 gnd
rlabel metal1 0 -299 95 -295 1 vdd
rlabel metal1 147 -337 147 -337 8 gnd
rlabel metal1 91 -300 148 -296 1 vdd
rlabel metal1 91 -340 148 -335 1 gnd
rlabel metal1 0 -394 36 -390 1 gnd
rlabel metal1 0 -353 36 -349 5 vdd
rlabel metal1 6 -377 17 -373 1 D
rlabel metal1 0 -394 95 -390 1 gnd
rlabel metal1 0 -353 95 -349 1 vdd
rlabel metal1 147 -391 147 -391 8 gnd
rlabel metal1 91 -354 148 -350 1 vdd
rlabel metal1 91 -394 148 -389 1 gnd
rlabel metal1 0 -448 36 -444 1 gnd
rlabel metal1 0 -407 36 -403 5 vdd
rlabel metal1 6 -431 17 -427 1 D
rlabel metal1 0 -448 95 -444 1 gnd
rlabel metal1 0 -407 95 -403 1 vdd
rlabel metal1 147 -445 147 -445 8 gnd
rlabel metal1 91 -408 148 -404 1 vdd
rlabel metal1 91 -448 148 -443 1 gnd
rlabel metal1 0 -502 36 -498 1 gnd
rlabel metal1 0 -461 36 -457 5 vdd
rlabel metal1 6 -485 17 -481 1 D
rlabel metal1 0 -502 95 -498 1 gnd
rlabel metal1 0 -461 95 -457 1 vdd
rlabel metal1 147 -499 147 -499 8 gnd
rlabel metal1 91 -462 148 -458 1 vdd
rlabel metal1 91 -502 148 -497 1 gnd
rlabel metal2 0 -240 4 -175 1 vdd
rlabel metal1 -9 -502 -5 4 3 gnd
rlabel metal1 251 -1176 255 -1166 1 A
rlabel metal2 282 587 305 594 1 P0
rlabel metal1 258 708 305 716 1 P0_bar
rlabel metal2 282 175 305 182 1 P1
rlabel metal1 258 296 305 304 1 P1_bar
rlabel metal1 259 -112 306 -104 1 P2_bar
rlabel metal2 283 -233 306 -226 1 P2
rlabel metal1 259 -515 306 -507 1 P3_bar
rlabel metal2 283 -636 306 -629 1 P3
rlabel metal1 90 -216 147 -211 1 gnd
rlabel metal1 146 -213 146 -213 8 gnd
rlabel metal1 259 -920 306 -912 1 P4_bar
rlabel metal1 374 -63 382 -59 1 P2
rlabel metal1 400 -70 409 -66 7 P1
rlabel metal1 371 -38 403 -34 5 vdd
rlabel metal1 371 -38 438 -34 5 vdd
rlabel metal1 371 -79 438 -75 1 gnd
rlabel metal1 393 -45 397 -34 1 vdd
rlabel metal1 374 -114 382 -110 1 P2
rlabel metal1 400 -121 409 -117 7 P1
rlabel metal1 393 -96 397 -85 1 vdd
rlabel metal1 374 -165 382 -161 1 P2
rlabel metal1 400 -172 409 -168 7 P1
rlabel metal1 393 -147 397 -136 1 vdd
rlabel metal1 379 -216 382 -212 1 P2
rlabel metal1 400 -223 409 -219 7 P1
rlabel metal1 393 -198 397 -187 1 vdd
rlabel metal1 374 -267 382 -263 1 P2
rlabel metal1 400 -274 409 -270 7 P1
rlabel metal1 393 -249 397 -238 1 vdd
rlabel metal1 428 -270 432 -255 1 G4
rlabel metal1 371 -283 438 -279 1 gnd
rlabel metal1 377 -242 438 -238 1 vdd
rlabel metal1 371 -232 438 -228 1 gnd
rlabel metal1 428 -216 441 -212 1 G3
rlabel metal1 377 -191 438 -187 1 vdd
rlabel metal1 413 -181 438 -176 1 gnd
rlabel metal1 428 -168 432 -153 1 G2
rlabel metal1 371 -181 438 -177 1 gnd
rlabel metal1 428 -117 432 -102 1 G1
rlabel metal1 381 -89 438 -85 1 vdd
rlabel metal1 428 -66 432 -51 1 G0
rlabel metal1 428 -114 441 -110 1 G1
rlabel metal1 428 -165 441 -161 1 G2
rlabel metal1 428 -267 441 -263 1 G4
rlabel metal1 5 17 12 21 1 A0_pre
rlabel metal1 5 -37 12 -33 1 A1_pre
rlabel metal1 5 -91 12 -87 1 A2_pre
rlabel metal1 5 -145 12 -141 1 A3_pre
rlabel metal1 5 -199 12 -195 1 A4_pre
rlabel metal1 6 -269 13 -265 1 B0_pre
rlabel metal1 6 -323 13 -319 1 B1_pre
rlabel metal1 6 -377 13 -373 1 B2_pre
rlabel metal1 6 -431 13 -427 1 B3_pre
rlabel metal1 6 -485 13 -481 1 B4_pre
rlabel metal1 137 16 154 20 1 A0
rlabel metal1 137 -38 161 -34 1 A1
rlabel metal1 137 -92 175 -88 1 A2
rlabel metal1 137 -146 160 -142 1 A3
rlabel metal1 137 -200 153 -196 1 A4
rlabel metal1 138 -270 151 -266 1 B0
rlabel metal1 138 -324 151 -320 1 B1
rlabel metal1 138 -378 151 -374 1 B2
rlabel metal1 138 -432 151 -428 1 B3
rlabel metal1 138 -486 155 -482 1 B4
rlabel metal1 364 -130 438 -126 1 gnd
rlabel metal1 377 -140 438 -136 1 vdd
rlabel metal2 18 47 23 861 1 vdd
rlabel metal2 0 0 0 0 1 gnd
rlabel metal1 258 693 262 700 1 vdd
rlabel metal1 258 803 262 810 1 vdd
rlabel metal1 257 593 261 600 1 vdd
rlabel metal1 258 483 262 490 1 vdd
rlabel metal1 258 391 262 398 1 vdd
rlabel metal1 258 281 262 288 1 vdd
rlabel metal1 257 181 261 188 1 vdd
rlabel metal1 258 71 262 78 1 vdd
rlabel metal1 259 -17 263 -10 1 vdd
rlabel metal1 259 -127 263 -120 1 vdd
rlabel metal1 258 -227 262 -220 1 vdd
rlabel metal1 259 -337 263 -330 1 vdd
rlabel metal1 259 -420 263 -413 1 vdd
rlabel space 260 -527 264 -520 1 vdd
rlabel metal1 258 -630 262 -623 1 vdd
rlabel metal1 259 -530 263 -523 1 vdd
rlabel metal1 259 -740 263 -733 1 vdd
rlabel metal1 259 -825 263 -818 1 vdd
rlabel metal1 259 -935 263 -928 1 vdd
rlabel metal1 258 -1035 262 -1028 1 vdd
rlabel metal1 259 -1145 263 -1138 1 vdd
rlabel metal1 196 -1053 200 -1039 1 gnd
rlabel metal1 185 733 202 737 1 gnd
rlabel metal2 179 360 184 670 1 vdd
rlabel metal1 201 585 220 589 1 gnd
rlabel metal1 185 321 201 325 1 gnd
rlabel metal1 195 173 203 177 1 gnd
rlabel metal1 186 -87 202 -83 1 gnd
rlabel metal1 196 -235 213 -231 1 gnd
rlabel metal1 186 -490 201 -486 1 gnd
rlabel metal1 196 -638 214 -634 1 gnd
rlabel metal1 189 -895 211 -891 1 gnd
rlabel metal1 196 -1043 221 -1039 1 gnd
rlabel metal1 364 -1187 368 -75 1 gnd
<< end >>
